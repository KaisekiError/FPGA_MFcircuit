--
--Written by GowinSynthesis
--Tool Version "V1.9.12 (64-bit)"
--Sat Nov  1 19:49:11 2025

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.12_x64/IDE/ipcore/FPADDSUB/data/FP_Add_Sub.v"
--file1 "\C:/Gowin/Gowin_V1.9.12_x64/IDE/ipcore/FPADDSUB/data/FP_Add_Sub_wrap.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
IipOOL5MTidF5RR3rDb2X7ylXa7qf+m1uPjsYjMtprPvdOxecO/b0M4M++BMT+uMHLvh88xytQ8y
rhWh2S6R8WOKehTgTnOSn74GLMXZ8NmafrhvpURKs8C3Nm64m7qZYYbYRJHz7+gOUB6cVrxmvL9E
0U97MIZj5wTMT73yQV8GRqxalFpTU0iOdXJXGyhZ1uQcziYD98Usnko8GKPo8JshXXq8VGj0UCsE
df6HY2hfbEgEpprKlV7j8nfdwU6gd0pTdXR9PLQVjjk4QNRG4/IL5VleCKJ6tbg9UnENU6CMXzqe
ZY/3JgWkPAHIMMFWGCvHjtSy2LGogC9mE/2WlA==

`protect encoding=(enctype="base64", line_length=76, bytes=309824)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
8YtbAvjDCysX3J4YlNajdVtOnhI9ZEmLBAwHdyX7g//4/Ur7rl5bZha7Q0cvZhzhCBMdXjeKP0Ar
nj/lNv8VuXQDDhtFfN9T0MNoOX0Wt9E+FxCH0aTMu6PKVv9kyVHSQg8zTl0+WxTpCbSdNAwkgjhQ
eeBARBSRFUC46FdvK4ZoGDac3INe5VWr1rdvPqMxJDQhaOelDspjsohjHkGg50wDoqcoxDd/cOrs
ou3sVpru/Ir7qgcg6q87di8quY53OB/BYEd/C53Q6jH7/Z4Yo8BdEALSZJvgY7hLoHLVQHBwHKXz
zJWhzgwH8bs2IdPVx5fG7bwCTBI7rrKfDD498pM/8juBy/5ixGsUk9Yq6IzMDRFzPlznbbw6ABhk
YaI62g8mZYu8SzRcH+d0PvlYWPQHKsWS4Qr9nGY5uSwREcdzKJKoYW6avwbcVEJwaV6qwa/TZU+7
29KLyy5oMpOc/aZxhxLi1F/WnQgoG/Ite6kSpN+6Titg4I1vc+5HlWWpNUgzHDnjCIDCTnNSzPBT
J5R9gKiXCOnb73NvKg+8j0R51d7e4D1Sw+d9rC4sqh3XbgY0DomkOhEzSN+neNQYyEsDTGmuW2Cc
Zo2rE/BfIYogs0eluWk3HkHXJA9uGxNAU5U0MMwnrEJTt8kYuBTrU8sLL3y1Q6q1+6nphs+d0to/
II8k6sC6DrMawtV/84yMnxpGdqj6XwhXMn+pcYhBFENYs9YvK5x7QZzaDxMD0Pk6+0w9jvrqjS/7
ncPSKuJhR8KKIoznevt3r1Lab+YhKFhmu3B6IbX/MK1MTRMoMv2ysMx/DCU/0oVWAUCYHT4kzXAH
j0PyR71a0tXZ/ByJIey73b87JLiHJTjtqQgd9uYP2uwb4VtOobNMlM+XAQuT3blhy+9eBUElKZ42
ZrXQw4bxAkXXRhxYZu6w10hoXaOadQhVzPB1aZ1ppCTeNQfmv6VkYFYMY2F7/U5ZrkfKRs1UPy2Y
6mCftPWYeUGFuGyxBknm6mrVPiyXC2wGuAyPG3Md+AJq/EA3M/p64XsFWABVocMJaPd5hYJgS8hn
SMbk1t0hnAeINFJck8kM/eWtgLZVCQJ1I9mxStdiR88qfu+j0XzNM2uc7gAnHFomzupRpxI6bJQ3
z+MeRTln+lzK1YIjspBRJ7hbZmpEUFd/wf1gA3q/YgnlvnskeNlIAhg6R+V1h+7IPYmrEIPMYVZE
cfQxY1R70Fe8M74ACP5hTEu4kBuCCHRHtZtN/wR2OG17MG2ODjsI4EBHy/olaY3+M0GXif1sk0eW
KBeWlxPdso/rv60E69URoVLTm/Fhep1/CD4I6GWRXzr7o2QOQHlLHEhIE3GNTmZLPNZic2mrD1k8
d4eLg4OvBiTAZJxwTM0FQcERIJiKJI9BNABtd/PXSxKyQ7KqVDOFUjvVFg8OXio4L6V8KMjSsBuc
xEVD6InGPilwoCHBuKoh0kvWi1qvNcHUUlNAoLLsdDxRIR68hXAJ3i3iZWSnznBB96MD+Mv1DiR1
i4UM8WLAKHRoaEwVelh3y66zxUtUSjmW2bjYIvhCNNQIrCGflU0oKEGaGfRZI1Ih8zBLYiZ0QYHN
qWvd2s8V7F9sw2SXCefajTkRFC+DE7z2pe4xes29x6Xlgndoho7eMIv0avVSGD9OfU9M/wV4dXc2
s05jZQ2d9u7OqNzyAm7EiwQ/4edgPL4joVtF8YnzKfoj3RX4u/MzIdZUxVUzzX4a8E4gBaixQ54e
R5AlXWt+uRzjDLZ+2O5gJZjHtjLAvzgEgWcJYca1nyiq/eOfN8gTw7/3E1SvldgYxEOPpm7s2+Oi
q+NxGK3jFaU0Gt+kzGksyyhHlKaNYiAS9aTPSM3GHHZ0nz7c6JXFHBb/sjUWz0DpeQ2tVYORnp4t
3MlfB4/k6xBRKo+DfPZ0gJ9JYkmWDBh5KUO9bsHHwRFHZIYIS80G+4xaGCUnFNbeKFDiHmIVKU5G
BVGioojQhIzEMKB/6cRWGeYehSd3kWlEXhYcQWZrLhK6FJ135JEWcFKy6SD0S6i+N1zPPO2d53+x
75WwkcbB+eoPbK99/ooBA2rmvGn8QncW/2jpxZiOkVuUza1de8Jj7nW7kMcXmSv3fvfu4OkCioVM
AX97wPKXE8JcpuSQiSXkm4mCGXD87tqPJIdwtC1hn6AGRAwCdP11LCUY5DcJpB0W6OXPAZFaAz+u
gA3nW6tkqMNZI95dSQnMcNR7xuNys8DKU+NXJZ4k26AY7nMsaMolhBQi43ARW/sex9EhLRH3yIng
NYZE8U+ssTKfS+pIxhoKu7+2Fb0iyNE7CUOSt3ZqU/C14Stpbt9pssXQmjiFNsKupa6FVX9k2uWQ
/CZHCZ6TopmoYT2pyvRCEkPYwNsjfht/WJI1gconZWJxkO6LhVkQq6cExY0ZY51OrF2kVZ9rwe27
D+SJPQe5Y8eVrRM1bIOisBseOagPJmCcFg5VqObhaaKtmZQYjtKXMchlfBoFHAOcHoFbyfcFWYbd
IKqgC0nXqDYSQ8zPb8LS1Uw71be3x5o1srxEpv/lLDM745VIp1kufZRWU8XcGz2aFWT5PRxa8xdD
/mBIsO0jKJCbBPXshxBGQlEY1/c1PMZ8qJTjTlTW8WOx561+MEMJaFVEpX44L1E2gIaIWKEbmZFr
g6OTio5J929o83M0mhGrQvAI/NVgwniqJe7DTQRqYMXlyx9rsDQyo+apAcAI3A62elFemOcWMh67
wXUdsXWFs7L2F5yyKpxQZ2szHSZJYEor3svDzkEUhAabgFCqXU8b6Yha0nldahKSD/uUv9PCyXMt
y7m8290zDvb9Ag50wcJX3DPUiDkS3uqmHv9p/co6leo1/SCPf2GAx7GSGRZrAMS/7tkuA39zac/C
dAw45Vh2Ht8ElhUGm8emPIPpR8NnwdjfRipJ/SexVUr6XXF+21qQnNjwEvm6WekPN79mN8n0feTe
Iu45+/EGSvI/8SP0cyo+6phLJ8PFSF9FYO03QXe3TyfK4CWHVADu7TCtp1gd93YNduK9W7u9xbZm
HvlpZeuc9iIxoWVwFabTGp9MdUs9/aacD8zMUxsYQmsCLP27h1tcBgGoVbHzC/PTal0C9MrpOR1Y
8NPfhclPQLbTEC332iJ5m7cf2JWbaxgGXAmfLHQCmHGY2bk97HbIqbHoLNH1JTWmCecnV6uE9FpE
0KMdX5cyUzUKirjJsrDlfuZfsAaeMK0T338d1ku0sKxUJ0cZHq9pc44SewGjbzUyUBPirOvH6oWi
cyMTrTdPCjZ2l01xDMO8hGpleRAujkb9vRO8bAhl6+KmJWBxLdohV2pIGNFHw9JRnsviQrES7+LF
kH05XnH9Lvmzk/DkKG4LtHX5OZ6dPYq+vHp6CIZoML0R6BJzm5OQfqrV1FsaZCqH8RBzSA63d46h
njPyL6FT0AfgNmpvP9Vc3eJ21teEuXNyie6TxlJoe4xIwnBPT3DhP4Ltc8ki4wRGcs46rNvtBgJ6
LyuYKdsav/FRworR8Md92y7fP/phgrWOKBcrddTpYunnuP6p8vmcdx6FfaxQG0sm8q4xFwzAsfx1
Sc8PayRbEWd92jOGUUDGRIAXqouRXtfr7txxAAuTZzMWc3tFLFt6pXiEugoFJwpeWAPoE5WEjtqF
XNJR1gYpYDj4ozBVkfuJpDYuKxXhAi/Zkv97yBapbid6vVn4pRj7OQrWFwjeHBr4llNXW6rjEhYD
gYZiS8lY+gP2DnfQD6wzXVVSloACSMCHv0lpSpHMEtGAgY1Q+GdPYnsDna1hvnH+fI96jw8n9qaC
vtcfOc3CcsX7zeJUYmK7cVloY6tZ/rMDHo/tV/shsrvD2ZKFt5ghv/QFHqCXijecirDEx7eKaTL8
AYUdvd2F8wBZPYm7TucagQUg91zn7xEoyIKji9jsdHDCdiaH2WGqn/7wl2qkFkUvESuFzMJfiz6S
V+1VE/5/wWAKxgLRItRm4k7EyH6qhQtmGj3WOLzzaD7P5ipyEf6ODM3Cqf15QCV6pfL2G05MP3JA
BPa8vxtUqUBTg7UXNsLDUZ3h3wM+vULAd0usncyB8xkkQUNfyj5Ij8qdczsZBWoI7U53Y/cyT/ta
eFpz9UqYf7ssAmGktujR6UidfbQu6u/O84ejo1ya0T0vBnVq7z2NFVMJFkpsFFKXDcTvwB5BOYql
Nqv8wCHoNFW204cEgRAdHusFprQLXOT/B6Gqxl0OmNaVuXy39SDc3um6oIHNAZ0bWsM+qGL6NwJB
GSXwmEm0qxpSWZHSkuUpnWCEJ7/XftVkpFuU/IUHYwEcmIFj/f0AxNgskp16e98yBvCU4dwacvCp
+5oaeLU1qNGhb+VK0bSgrOfTkQQjnlRrz/bMCpZH1H7cVTj1MkiSxcBYbiA0BLlxFtXpiLDDIYon
VmgTxzHMONyun0u8UXAQa/7VQ+ZfCC5lJ6O1hMBhplAaqST2uCEPRwF362/hBOB4lJD/JuDFznwy
9THLxtGXuXZDYe4JL50lMn6a4sQmqLkl/kftMH7ZtJjVY4sMgOs6qrjEwYDa1q1PvzKPcKUMk4qY
OlIHAJpR6xPJ5UkDEFjZ0zZ0aRn4FYtw3EsZvMxbKh0+L+qmrSdfd0NOLG9mkirAvVGdCvSNF4bd
eWCAcycw3/jKv2k+KidkWEIIuJbyt9UGzsd9UPNiqmsOiF6kbDquzVxfJPoQXQX4uroU5zmLblEj
zS4YGtWN3MiUCiNISn2laZP0TjA/5JtHNY/UP2ruJSoSGbt2e2o4QHi8X33VHdb69NfXzwCdmri6
UlPj34OrUzqVQrENaZ1jSXX8wdHPLc+CrZ2Xzd3JffLo3P9igC+7ZwYKMcOn+nMvUBbyBQYe2r5Q
2Na/wWRAfqBFSEGmkVOCz5faBH8jIXnS0dfsduv9PzvsQ4YT7HdQ3Dz3sVhwdrF2tSEBqakD4Z6y
r6jXnWQxAms4GmU5hcr/dUg5pybiPA6rgJ4gDD/ex/7CpW+/EHtuHU9TT9XtvdApxTdu1EQ2hQiv
QYDXg4AHN0PGvUQrSPtYMpevWhNnqu6HsV+5qfW8sLkhfpMNJ1wE8CNEywEgcJJq0x8UcKw4CYf7
qCwqJOpRPBRP7GArHmqDX/Bvjjy7GFwjBCDzN65+pJHKHgp77PlWKl477Wuo82vWl2RnvYMpjpOY
6KTqEcCS73SGy8kKp12xusmU/iak8RbjCHu96loFWRjJFjtjhHX2C+/HTYHGyAMGryMIt1SyDkL4
aKTWuPYcuIXURnyc7ryuTJ30ymitj7/ukXv14ecvHSN/4ZS7YTA5hhkNAF9ms4YO7TUve+q7ma73
INyuSofAUfQ0wdIz/LxhPIy3v0rrKRtdl7654luZj4g42aQkqGGppHlysVE+fKgtdN0Q96aFkcrL
dDTcfP/xYU5TLTeb7+87/GpL0kin1SeehqC48WwayvbYmDtdmZy6/Ch+weWo0lPo43dUwLbUIahD
CGYpQg3GSFLlEGdZuqyHSwliVFmtVoi8O3nQcHZX0rv6v6wQB/U9WdTH15LfvR6bX1ONe00sXdGQ
7bZdXu92Snwnh0zjRCIZJBEJU0DlyaCEKL9Et2nRvpZRdrLfktYqwAI4JMAeLtNZbrjVs3TL7yTF
22PpAzGY8wUBZN1GgbNQF40z9ztEVt5S7asD2AAokEkVKDW6BPI6A0RXEFktr0XSB3j2/CndRBp7
55lBlcJTKdrlBfWaxWf1eStQtGWsPsO4MGgg6H4Ev2MIiW4A2GmlZlEP2fFvMRkFy3bOq6MA7WAn
MgIt0nv1CJ4jI2Dyk6cp2KW3q99CRn5NS0eruqK9I6ny4j7WWxUrgGLCkbsbovy5VEOox2DDvI5L
Xa8zqjPpgRQQZaeAjTWJiz114hjiou0juKLnUTi2218gbhaurKes2G5rSdVC1Z+v9McN11cw8ALq
qn0Bq2UOvK/vdIho0LM8fYh4pOcgrVcwKfl4dXXOEK02OnvdbRzL6u08hwlQKR5FgGB0VU0tz0bd
l16I/oezaGq6iYgtrWiacmXkzG3wifHG2gv3GsInQqetxjFjp9eery0C9zsMGm5PmNnaKoYeIqUo
PXE+XeMmsEccl1ltkHATeUpEnVMyUD3YGeX9MCy7swmifD5NP+VCkkkkuv4I51OFqv+zu7PAMjTG
qy5gLy2USFUKJ+JXOrKP8vCc4bvrZ1zjUMW/NNIEf/ztO/K6gcw+k0mJAinIgxB31YyMYSIT49C8
q8nz7Qze6IW7pzabGMr4/CqQLYP4rFuzlNpuYoEfF1PPxx7LbEzxmMLsES8FqFXCZpzL77BAG21b
/3XkREEPqm5YQfabVqBjucWRm74LjMjXfH00Y6vOapfRR2lMOBWeU6NIx/KDZIlBFRQ3ZI42KOup
5W4emw9KJmid8WXhd08d40fiDZ5ZHbUdTVKML3N4OU4MXqnHcmzqtOTxNOhqy9CKw2LxtaQoktn+
Z+eSBBKtMBkSf0ir3wFul4GGwePY6y7cm6+jfj4Vj2PheWpgezaBaYG1LRBp5Mr8FfPXlTiKUa7P
QKg2Kl/VUuvS8X2t5lgHtTXPlKq7xw3HWdI1pZgpIdurgorrcLQpZtnS05RdoLPGy8XyTo4tbr+6
512w6fiUc43HQnQSK1Qvlq+8/dRuLYksVEKCGLn2j1DpMB3cWkvHTeYUnlmOT/aVv1lZ++FSXTCC
7qV7u9HgywZ9hoK8XLINsL5GFaUH9EISwPiQjYHV/d5DKknJgnfaUYLankL9m+ETF9nu37dvtY8C
Mx++73jEA4ILQXrLW3wCR2DGrxZnsQYP3F6g8w0fgOvymUpyW3uaZwjadnSQJy8jeHJgp7c640hM
kp09YL9Al+YxxskJz64GcRKJD7UDRkECzmxJKmabVNCOvqwfDQQaj1SrtbPngtIKD2Y3YvcB9R7O
9kxQt8A5SZlEq+XxL9rB/P8L7xUCOdYCwAHgb78PzrQDLUY0cf1y+VeGj9yr2vS2dpvH9MUsiBZE
vLQ5mlTc168yZfGrjkEZSj5xsEyQ8GGZDmPGPecJNw+zp9dnDaUMZGqGqXH7f0/tq0RiaLXQArbv
FvbJ+zhsbvCTV/yJ0EONdni/vFoOFJnJjIHxA0sOW7bJvK13lfVGRxTFCQob6pmy88DKVCNEScVj
mGI7i4X3Nd1qLgkrHXa+SWuBBLDlxdSKIpnsfkMQ1+RiNzZvyZNsXE3iYb7FDPvnW8WFgws2Y9ku
woGz3lHw2xMU/PqwUAQml9xdMFVjXHjJ7HUlIor7LDzhNcg41f8gxEDPsjC3tFSjdqy6Q6MjFts+
LGWe4CRT3pRfOjPnjk7/RmNCLeBctf5N2QcWBUFHGwtO3MQvbZOUYB5qtAqkiBLnrovimmAx7tlS
LWNsQXkHQX3RHYkpXieZb54BWdfoK73xXI2jNSph+5Nr4t/E5SQ9OHLARzVOUqLjgpKp9DD8YVXv
GPzmqvSt7snij1dzJCWb+/1Z4aM7a6c6YBLiVaILSNNZmbJ3w04oAp94COw5nnQRYW6mBDboEqXQ
gWaicXgDVZ4ermbOptF/MP9/sVG88WqL2k0jAgXyjs/PQ5cepy5hmUeW08KrzRp7D+iPg8R3bDkq
T2pfPqrNv+cJtlPDmzwrHgt7DUMR7wnBuDVmAGf14sz0TlREBwbClfsmmUTHsd7yq/lBRGGUk4b1
zO3WZ+fw7atNbJQearFL1MIQUcnI4wP3cwUVmwOiM3kdCmt6muL1rCUJHOp0lyMTp+58Uk2wPLdc
zamEPkaD347Ingg8xUJ/es6jOeEIo6wQHtBzTnLkUty6dzZ6SOLxq/5XU54YhX1cS6FYPbRecVvx
YUYq+wtMlWisj7+SY2qqHae56WisYR8vk0Mho5nAyfb9Ku7rqbiG284lR65U0qaroQlYyMsEO0H9
a+/P5VcsVeT9ydy5uwIORakgz5XCJx5bLaXGgh1A3q//X8LVn45FwAKEr8HcfdDcxOUXhE1whnEf
LHTkf4F9HGwUGqyNHpVI1MefHOMjHQTu+NLDrphFSvmtzBg7/AwdothiW8MSbSh25w7trCDekDy2
sSechtwNmr0vA33sfGoVPXcnoLOged7UO01I1aHdbEN8WwtlCwEqYRoQlgVRxjrs3r3MvrgF3/FL
IverriUSrgXE07I+xJMT+W2QJyykK+511YIoKFb+QUqlCRfKBRY8KXBan7rJWksjl+JlOa/CmwQY
larE74l2Yw9x1FTVzBehiQl+fO8jMpHbaP1nougjuTScNw0zkSzpWNVIdCJ7y28kPRJ1NXk40+F/
CzRE6Xd7gV3bpy/nHP3Z6eoyyVOvvItQyYegoi0MQVLltZZg4oYoAu5CNMgmw7QaX9b5scbYBGxb
qenNPbzjlL4m2uWiSejSkSHIc5NfvSLB0PCE0WDED6s9e9nwJctErvB6PDqoar+T2JTOWmkr/eTD
9ajWTx3G+ki67eM6XFWdiHiUW7l4tdcRzW/YO91oKHrKbeOmKUKmu1SPgC/YRfLMRi6PWaGtNfNJ
sqoJFZ9oMkOcs4D3fasgvkshel2lGJ/HTkXMc3L5XshO0U4B4vM7uvR4HsXMm9Tm9V5vRG7T+UCD
bQOGe68xaUgjnSKiedoAhsKPpWj93EFMeqLGXJAd7TdoL6r2U2lgE1lFVhIR4Ch3EKQu7kjema54
fIWoAYoUhnJUE3l9/Tecqg8OfDalLRpSdRtfbPOQFXV9TkxRV2Ierm/n7kBnh9qWGTQv1Jkl7AhN
MYvhCSGWLPflZeMiCYO9I0KYND5Kceg2tL7wEAv0yUnkhixpHEBli+A0LfuBlbvxweeWgwXkulpo
wygymB/rB/Sg4cPc4aqx47j5fzX0N1gJ06v4wfyY2nhizvM9Rp3CleDP9NOg10EVwQ+5ojfzicCS
O5rBQ5jT1xOVVJA/DbWOzcxKiyVlcCavLjeH1b40s1IItC2gfWQn3/yosbv47Cvcl7z1zjxMP9pY
K0eH9ATGlFUcx5uKCaTGXPD/kX3UyK3dx6gBaqMJi7z0LpAjmoMlSjNqNYgk7gHJDiuxZnGm4fhs
vuJfc2P2TwLBI5PEwVKSl3KzxB4XAlRq5PDSARRiBY/G0Pn0M3l4XarnH3y8N5QTklVIGNCpPY9e
8/6VFKEPqgmN2KSgJ24mybFIEfLpiYbTq2FDkRFjy9zGu42J0p9p11GSxaufe8rZerUR98ftsyIK
4CQF7pAICOnnqKf3p8sjUHJ3vMueTg4OGVt8Qtbh+PsrKFvvpow5De4gehstbHPWG7spn4y4B5Bu
DpweSXlC5zwmWlQe3BfpyLm6P/9z5gCVf4X3s14d+OUlqI1r7n0ywXDWIf4RtlQFFVYwiDBJTUJW
XrD2kvF6HplG5C35nPUNQWRVTFKLmlWZ2sUTmMexGlAb+Zw4dtnwefUIT72kdOmm0Q8N0aGXpGLk
TKyoRY2Ch1YWP366lUyTedEVtE/OunJMkuN8RhZl8jGcwBz1Ia28vdh7J553iIBPRyDvYhLf8Lx5
MUnYqPpKZeEPlUkh6poG5hyw05e4eRpmoVfAhHb/GUGew7LqZLTgBNsRvb93UbfS9yOI8x3plqOx
2JCT2gWrkrhx1nOkGG1xznAWI9W7I/KDK4qZFDe3WekZBshYDu/cir/ynMtdPQoSrXt+L9ChHp+c
qCBKeb0lUAp6bha0mlYP/f8oKhCVIN+ZiwzHPlNO2uqfGCU4BHc2nNtia6viKspdHJvf/pn/rFAL
/hZOr4ORfeEdbNkEehoCvcCnelHOL1ZEFwyqmVEk8+YRfMbYqK1aj5y0ztm9uXzbaqNx9sbi9NFz
S8UXZay6tfA2OmIlYrG79Zopt+f9CbpboAB+Kf/axdShOJDfxAcYf7n9fxXC+Hq+xkq9Ps21eOLT
0E7uGFEYaeDUO7dow+lz0ikCm2u5lK2NCPndo2EZtvJOH0NgsZz20FVhDDtOmgFJV3hOd8QNbH+Z
GMMmuJ00LemOIJnQlYPN27qiJ4Ihq9La8Bx5+yatDgDI/uAzl02/Hw6tS+euLxDnuPyG/2V7ijyR
+FAyo7K54/sBi76D87KZm2iYfsBgo/DIIXUYmDNNGUFsnar/mtFK0njfbUo0LaeJGpn+rx6yeIBo
sxXuwwUPNFLJYhuGw+Gl5xHaP4cJLpBIKpsiiNV+zSeJemmm20z/5Z+wruV4Fv7XctzVrHW9M8m7
Qx3IteeuDcnAoBrO4tZ1hsBCmzrsTkaFW6YF6YjP9ESHEY4HyR/UFMLhinMEz812LbqBG7KGCYre
B1XWXrnIftW9gxsvd/mhf94S0PytaPy/LEsQQjig2i2kRAfKSjdCglsKOhzuR4U9cQt8/vtpco4h
9a98VItqCIvXBgwwZa/whwu8VbLFu76FldbFgbCX2WRxe1r8yeeMJ0bUx/jmjxdlbgzQlphz5abm
tfOT8Sm9BbaEbCixIXzr3HRK7mi0dEsvzQ5PZRyycIAkQynAh0XHwNveCP3NQEhgddPHQ0UQ2RDa
Nyly+GDkzKxu6AVaPoM5ve+6cY0loBtRQfHsvNoBNS/23REolwxSYj8sy+KzVBodAvwuAB4K8Xw9
GBZw7lXexe/H6cBLJKQzHDUXbyvDVm4CnZfU+wgRfungWrckyv6B0VEYuIxSu+XK26yIzT8WxYg0
/7Jj9bsDI+aVNto0Qh4OdgIjcrmZMyRYzABnvfuYUPab19tGUfof4TEGiIfqyeOCSHhfY0otyCao
mkqvjUsCLjWbhiUGpF5ZXekqj/L2TLua6KcBHmqhQzTbwKz1uz98g+2W81Ko7XJ2ecSbRD7iTEcc
l2GaiL44e88p554f9JKoTE5awryolS8hF2KHI7sDK5yDF9k+ixd9djFiaSu3bHzmN26hkKRrY8t7
dF3Lbu4RvAeBc/ZWEeG24gBIwkBw6cekxwwbWgysMhMd3rqd9yiHuzIyGsozH4C5mVdtCyROr1zY
HwH5xhfc4WtbLzA0TjjkhUKt3S2pkTixZyqaBRvqAnHbvCg8ocJgLi+taqi+LzJ1CI41rRt/U3Ts
h6jPOxtMK/7EXM76Izw/sXgo4Tzr/4DXBoi/MtFGicnNiXHCAJAHnsUPKqAnY3UriS3fem5py3vn
kKCj1RoqZF6dKpXU3e54yziSa+JNUrZsJxr98KSNJ8Qz2WyBBXfqtiI+vRW7tGq3eDjludAHToGe
k7dL8xFQ7PjKGhEJ1MWLPS61HiTn88JO75yOd6RJkFElYP7G/SutgNThEz7uYwpzG5uI2X2BpCpa
/HT4h59j/vs7GaT//arDlwExX2jw71kWVVd9RBgjXP7wwaV78HcRNslMvpCD1dhnvONSEb92/zwp
5HucPI1M1dmsAsimjd79H51N/6ctfQ0DpHjmxgAUWnHV6oCX7vTZQedDFEFn/5KPCTgRjcXuiFV2
9oi9hEXfmO2ovPP1JZdpApJucnVg+jKTi2ZCa8AEKi/AIYSuIHD7zAX7OJ9U9pCCAQmagIToFg/O
dJvB/uhaPexBvKTQmphkf0pHbMfLVtlzXgES+aLoBUnXFvWE6TV4WMCxncY8w6Oe9c7+R8P4bAB7
OQRDaUvli/GR8fRvezCvhHlvY+OTKNUStRtgFOrW8O98/+/6UjcBVMrAYMPgO+0jWH6OUiYIFKyA
ml/Nneks1jlgtPKmceZ+yfKqmoa9Nurn8BPvhKfuOjRG2IAY9iUIed8ZAAqhoWE/tgsj9sRasrBe
zeQb0lZ9GOwKRjOqYL2b30iEMhvFMDywn3oXv4AEoQ9gWtJdYphiejjdNWYGrQiOPfyJpEp0gPPP
tEyrMPi0UiLmlxBr7g5ZgeSt+XupzW2ZWeXDx0m/WmzbhTLXf5v3vEdygKVxU3mNCwDoBpHVUoV2
7fww+jliJfkI4Z+BcuWhzF7NuOuWoQ1ma7TkCSXlryuF4rNFBcaHSiiybTO+8xUjXAJ/gZEr0Hyr
p+gQmMM8XDueU+P1Gjt3IsI9BVgalrgXSB7v657UQHXFtdVpyWPOSu3vVzSJ9cVEEgEDB8g0Z58e
Rqc33NoEEcC1rVBFc3XOuRQIBMUSLOUAwFirXfjx/ugEReX5x7EIbOBfQFLTISfgKbpPAh0tvGRP
RHwiz4IMQhgfw6G2TMy5l3KeSQeUop/0jdKMJyo+mgmUh8pBoNzaM1mmw5NzrqwCRM6iyjuDDrGj
prd68UXayw6NhMuohW9+w1QBkP/MZbLbGWRgFSDN/2yySazmhug8Bw3TWGk/RiDIM6aImAeAgRVI
BLL6VptG8+cG54kklGB0OomP0W2X6SvUXFicOLGvmXq8T7NbpVlfINKosLos3SLaUfjmL4osFZG3
aj0jPLpaGudYTYHEv4HCszNsp2mOy810ci1D/h0aPp88s6k2AgWttuI53MzvvuQeug3ZswUBe9H7
f1NoBxAmhjdUAcdtMjjY4WbXa8+v0fzk9SvDN+JcqvU4FtoN0zUesO3g5S0ClKP8NjAdBzcAqaV+
4Eiria7qZLZIKsDg9Xy5Ddk+FCPm0GBwCt5cakvxxjfkYqPjcDhF2JPXBmvdNhMKm/OkGMHuwj0y
04NR4S6zOXTYwUGpAAGQiE2eX8OcncYdlHXE0t6VTP1be41QtRDyBMp7cPTWTWFPG18pSLrcJsSi
C7vxJRKvRqZlJ9msrBAr9GPvGW5Vgi7ROrCjMFl83H3QiJ7qB7ekGX+AAFqUkij7R0Ac2uJ+jb8Z
4RishsmQZdyKMtDHbd9eA2qTn3bn4WL15WQpxplpPyzW8RPeYcehAfbIUut/Ffl8AIWGUJh3OA2U
bDgyWOnWYchYSk8KE/vHFf5JpeVcJzo60RCe5IsSWmWURHPCfxqrIfUQCRLDH6j92Oz64qO2tqU8
NFeQKYieKFalBisdT6w6rXY+XLzI+3IPaVQz7aHppzAkamUT/kfDtDWN8NF2WoUWMyeuscCY3EN9
4ytHzyHK+sjhYYxsAtvJyAUpCdil0EWIbF8LRBAp/yQ4rsv7BV9xNDK+733zppNVgTx8ZQsa6RAH
t/CgkxBTJxE++/9G1qjkbfLp2jBMkrARBFaoP1YrDFBGz4C0GmyqT1pCnnVDkGI7veGDeY3+fPzo
+a0947vt3+2IhEgYADSbG8ghhQVQdBZgK9vga6liM1h4XJ1Tk/WK513W1CpZhERAFvgT4CTFS2YG
b8nKlLGiL+deZEUEFHyGlKZrACfoTu8qSQAw/84zC6JpxTP3Fm/2cWxWtcE+MYobNE/FPNMKLrzZ
0cFxwdEK51zJvWOMe/hC7p5i7J0WqHPdTXIrPJ0OXad9J1UDcOwkv63Fri1QUxjV2YfgFO8TWCsM
kkcCNV8r4IPigamK2Xbm6YVBlPYcXsgzxPs/+Pi9lnoPScO3msbYppYygqXYV5R1ykyjgFPE3yRM
YIxo+f8rEMebb2Qemm3WQjM1Y6ORonUbiUcp1hNm8/Ml172Lxa0IoezTX8ItQCM624UWYJQqAXds
QB7FI/+dUFxPN2WzxlXIU8igxV+Tx/PA5rsHxvW/c/Az0IcXgmMVzfqXpXCj8Hx5+bXnKXrsRcsL
xNPVAXVBmOBKuqwoadnC2UDJBVqPOTjBOb5XtM0l7XNcEYfkUhGByRA9QmVYW6y9ekjS6yVZsMfW
Fd3tL0CvKI21avr3a8aGM43B6D6WisqV8GxzBKNTdh9jtmasPLFmnhWHI/fApqaLr5yuv7o3hcbw
B4ErRCIyP2O7zr2tncWUImrSm1fYl8GqF3R3+xJLcZ+3b88BAMNGOxmUGs1CPTTizlN0tcmbic9T
B2tXgb/Nk9TAggdG2p/UQX1Kvq8zT9frYigDDe0WWvjGrFoGAqzW6PQGaS6XDuKNtPZOfhKWG2XG
FJrH/FsIxg5KttLQKSyLYE99ta7i4j/vsa1dSfLCVN5YFLgQyq19DxaIjPkQstxlN584Sx9CD7Oe
0DUwQGIPurKkvyLWIZ9RnOO3lWXZYx0O6PUcTtld2OnWOluACIvljIliTqR8Jg9dcKz/WU6LN83R
DL52KIL1EvUo7BQN0Nb5pMfVbGeW8/9fToGNrnugCyUxfa0Ip6KxfrkxTmeEVyb2A8QNxKHwGuip
nSMOY0oAn6I+JSBB57bSMvnzHPO3OXj9Rgob9+RI2SMsovd7yEO3GP4F5eAc1EcUNcmcrU/1nlne
0LhRoWJ+8jPdyzddPyi4Dod03/RvkjHiTs/e7wFjS8GgI+4cXcJw9D4YL2LrYaYyTOYP95B1l0Zf
YCasH6n+PLDzRWRT2eGWgBuOpn8pow1BMes94hk36UDFx1wXa7sjN8zkHkesUSzTSMzKXZvKa4gZ
UrbMbl9CR5EtWjANTcyhJd88vK1kwefHvP7m+lGXPhOARDIYYG47vttavVqwALeDdaOAXx6qw5mR
W9G1WKLpCWygBNBMos+Sryv7GuW0akw0PInrVIxf2lPxuywYrUYq3VpsaqwmhiWQ7gayTeBmJEnC
XposGQWgzVvGGFjovmZJWQoQ9jK/dhIcQZCCY+rCIhJGV682jTpvfCaC6Qn9Wobf4DNtt808BsH1
HjN57GsZ0d2VKhsknB37k9O5mNp/t1uq2oxfSm2QPfqvk6xyspK+5IBF575aJwJPe5x7Yn2WHwuh
+lU7LzZUt1/79SQHGUw2JHydAMWCI7pQMbdE6ysUuU+LjHy8xgJSjVJs9fHvmdUSBGlhr/467OyL
pJkZpyaFxdUyMwOXaX+65H6ZjxzFulPHRrOW+O9QU1PVUhDmKXLgwS6nNsHY41OFbQLiOed9lOyy
FrbcfofRo3koJBrd/0d2MrRD31Bs7Fs/qYofePd8MzflrfIjfF8YcssB2bhET4NCdbUjdCxSmxJ9
lTGOM0tqGwuWbVLK2hT0U32Bf/9L1m61PfgT4/4hrF1PPPM+uLQXr+5wgRece9TaH8KvFFTWuD9Z
UuN6Lhrm/fcjPs3ChZOT+kOrOvckrhI2sbeQZA4xqfh4+erwYQuWkVtkNA2uaGyEPAV5POiPQqAq
0L/rPSY1sTVwCHzZ0yNJgePH+Mm/Q+bf4rCJAWWikjGHpBr4vwXIp8O+VgNIJSa9gLjxYZtPNXGy
IsYWzg2/2lm/VolC2prUdmKBkbRC1ECRJK6FMk/8biJlzpxZVWRs+HoEhUU5Ic6jtM1qZthypvhh
LqV1IWeB9AWaa7p3LGre4W71ROPYGgxcTzgCpBmqSv6/CLDTBEIiTFHMT6GBxdEqZ5OhWuvu7BxN
UZ2Fdy/KP7TUxebJxDsPe6oCyQX84gTl2+/zhr5oRm4rKyaVdI9AepKZIjR6NdSi1JQm9Npb/qRq
Ag1GJGsI1WmN/Yiw5lIb47vsfFpYbJfOZjNHDmhMSxEOkewqWTP/GGezDuz6fJkBue9FNhFC4Bcz
/4F8yJP7o30lhAhF6XKJ5yD1OEHDcPrjAO3odue9OqhG5oWJFTsNjzJyg7zL4J0vyA9LkBDPUfg9
IeJThdHlFqKPr4PMGrwrvOneWpz0tf4MeK1CSOhtnZvtSgqkqAXIRkwF+qfgJ3LR7QGurj26MgvC
W4qeFtEZeE7X1DQ6RF5oCvvxFNtm7OYw9fDFbEN2AXDl2HKUQjhBP5uXHTlmfACbiF83vn7xFRfU
siNPjPDqOfoq1jZqh0Sahr9WxBEXbqEPEJ3o26Wuj8wOSAtvKy1RBJS4mvcKt8HvCAbIsP1C+NEf
SViIwV3VNT8kQLADHNbxkZBPJQHYnJqVJFb4WMKZ8xy70480Vl0+e6KbFfGF47id2BXAmcCaicK4
3BGx23gLYqw8Q75PgV2it4kOjV8R705z6K4JzIb+8hEYMSrVepM+ub8BV/bIt6WNu1Mf6AnTRHy7
a6HnQM4or8zeBwZLFGU8K3MIxvrsEA5FF17seXhGMcPAcVbJj8/qIbyeUpNWLWMzhGq0mRM9Y+gQ
vC9phQU9WKMq1n1orV90IQKNcV5fnXERdOHrKNr/tsrRl8Z1vv5KC+1n3VdrRJ6yhCMpcVMWW15R
Rxw550maEzqJRH/42+mWwELLN+GZEVxHJrXh+DhVNP9wqExx7Ryumu8m7igzIWE9YMl8ON5OavV8
07WitVbE+ePf89frItBkxGBDnWoNb52YQ1KLpVV3IVK3a28qv7xQPvaq+S6Ku43O7QK+HWOI2rtb
bEdG3t8JYkhGqjo+nCxaNENeKkhzVv+nXSdE58Gbw868IYjW72o2RIfg4vXfKc3nHKA/O+jJmBtO
6F7R7B1I/i4ZZjI+zdgIKjXMa9ZLi/rIVqfDkIp9A9gZ6DTyO0iGr9QVOZ4048f/V140Sgn367lP
snv9XYgE22+vzl9xn2/uWzU0l82Pzry0t3wQm25qdAN/5hOT/vnuKLSFZyJasfyF/g2FWI9XwdKB
ybvqgJMwB6OL+LaOD6WhzEb3ffNHDVeVSrT5yDB1pzlr+xGf8HhpwUkuDfzjeNViSzz/5cdZHEDd
otJ1Tee6TOTJP9ApPQPFh+XYTuqLCm1RKaQeIIFBYBGxFNK9dEplklfKRdKBHhyiqQh4Hxitjw4l
X1Uazj3o9D9PpAlsDQ73zy9x/bLs41HjNjUKHjC0rZt7lDX9vfuPv2oSOYy8843LgQCYf6qEscG9
PWayPBXC9cJLHIqzPQc4Wx5VBscGJ8XOXkfdF3fNonwPADILnbS6WS/oPlTwpnC27Hcp7kWtcofp
gKRMvYyKoUhYxsGtldd/EWeFtr8Y1CVExjdfrUt0rocqH2oWDXOF8l87++qJ2Oqblz7Z/ZLTyxS3
fWrMxhzCQtyQf8JpyjdrgI0sUM2dE5IMmFZU8fbRw2QZy1lJbfsUt90LaaIANZc9ez8iq1a1xrS+
tS8l/KAJbyuEnB3KtzGrcciPBMDnkPvz+KSYbpwxtOiHC4dd1K0JtjYLaCbR136QzxLdCiwWcgW3
nQMUltjxr6dRq9TRPnsoUB/MPHDJ/y0RSORoZCM2WWSSsI5mD9qYfcNe15//S56G0MMa1ahwfl1T
Cantj8IuqHfycX6DJ8HJw8koTu4I30m7vs/H61QEjoGzwtrvB6rt21tAo9Qa0rHtb+ggToJc7UbX
GtuPpCaJvWDzyClKlvcN8U/0bPBeWda+HJae2e5Icw4+/dR1Jejo6NRGfTHCNqb3ehi6D/ww5Rrr
TXqJkVYNVBvOHmR8rKXX2mf2OwxFUWoJe3l4TREM3U1f5phLS3shBjw+fF7fHKKtt3HPtIosI9HQ
bH7wgZumGYY7r9Q86rGbJ9jF28SS/HB469Cf2t5JM+BDzK11ndDMTKHIZBg8QPM3vG24jhJn0Aq+
a4n9v5nz1BvxtxCncV4rfk+9LiTY0uHf65Ps3CeqNnP8VayRTuvf2pImM+nUCjfVNdoHTnQ+qb0i
Qmopc5fjUu90yhHjS+OawsJvfgWwIM4yUosbf+6l8Wa1UW+MITqbVRxdVjFJDywO+JBxgPPcDziq
ERm6iTduoobZDCTfJgAdL59Hhx+rLTunnzD4SaF5U8nkxqsW2EPXB9jDN24RdMiILOutk2UHu0YI
pDj4bw1PjKVQvUegpWvbHjHfFuZPJ5hrqfYollOSDNhyI5a3CQ34WY5SxdUYS/4JMd0xrkTxJrdR
Uj0eQk+hZQnlCttAJHfPqCjG1LrDOZH3hCNI8v+U2fSnNfqyvvtm0BML0fzt+ybYloWDxjuEaK93
IWYissK6/7fHzn2UxEiFbdLzaAwCV5ITU2oifwh5u5I4emHoEkPfpQyE/kjIeC2JXPQ4ZDEcCbv2
G7mGIe/gU3InJjZtDZSskJ6flvqkudOPf4J4pR8N33jNi5qNaazjzGBi9Gni4HUOyCA9UPINObZU
VAOV/KkdD4JKKTxXRLcEPyhELK1nAxnBZBYlbnR3ZqBkIgmqNUKFn58okKBMkpoXQ6x97JAmPrUv
LNkZn4ixbDa4IeULQSTYnXmn7u7WIxc02A9s+Wsrm/4xoYj1Gaxl9/4NU4las0BrOUFP/EKvMZNn
4873MDtUExnsL9oNAc0aUqipFcrozuhjRZK2bdLeq3endwVxA7R0t34JWa8Rzv7S0Jsoz1llzK3t
PcDB3NX46hPIH/2dzeOZpwku9YV7jhUxFT1m9fRmmgTMQ6ME4uX5MHeN9snrioteHHw5ZAxLrb9y
+69nABpkzWZpv5Ja6NsBTXKW0qCMsEvgairMTSOfusMbuICuPrQzGnyKWAo3naR3MPLUnG0Z3wNv
7i1h4gYbILnJZuv4/4aG+1NF147vkLN8Dejlobo8nNHJo3ZsTUEu6nJ50/K/4ezb+RZ74RwGvblR
EfngoM+bbGeiyN7tBu55XtS2ZZ+QENuajXMPhyl4L13HgdeYfszf6yYlYtT7l8345xuhhEAjyDgW
qjl5OsfyOXaR/f6r+VVuFzXdrxDiX9uk2h3CbixDbbAnEc7xsWmuP7ZaXP7/KUwVj1cRfZ84vmZ7
RMlnjyRO4YMuJqJeV0DdfnqnI9ljW8X1UPURMo8N9wzMVfKvd48RIlo6FKjGQKMq2RS0OgTv4lJY
VK4odDgEG8WTmku+/g1VG6Pyts/F61rjKDj6kRDwRdlPWDlCr0M+pkj6YY/b4cLTTSdZ9l0Q3K0G
p7BFr8xwwNjAgeukkB3/ImlC/QcxKoMGS4acJujEl/9JEyyIQK01bQRgFL8y9du6IuKbjbOTkxF+
eRX8nWgcvqhhFjAr4qRgOwfrGehaiPWlfxSPzrwiA6yoP3z+dzE+CVhN78vwVQI6k/02gseoqYQx
ojCmQXsPJSNrAIwrYkQ79OvR30EtcA7/JtqPL7BIDwI+uWmMpLjj0O8zAL6bKuKed7WP4UQemQyw
9oRK52O+M451VIl13hVFRfzMybjheWJ7CEUG9Bkyc8Z0R8LJqTbsu1kiZXgf/yb0gf/l405Cw8Lx
3TFCRBW3JBkEUmhZSbXqJQXQ1wWCOcYjrVVZmJvZ9ChHOTNbujStWzFoJ0pAsaqh2fCwh1N58Jkt
NQkkG9ccvty35wGW+rkdDZPhAiBKvlLLgYR1ediKpdDpcvhqTHuMezLN2SDkcYTjX1/4Rp1M/rAG
Kka7sMtJDv8N1ubBo8eH36buz7+fDd81BqE+W4R7O2/I223oCM7s1trxVbR79bc8MVHi4Ju9t3R3
SHcU4k9StB+uYjC4SzPF1uB9LdAZdqOg/nyoAnB9N0rZfRU6BJjhTT1UadqdoQJy9E7Vz6PcY0sx
Oy4GkVis9PpPm32TVmQVtdPsIy9AuY2rYEA1MISrm06sWxRCuIMisg+k1sCGxr6FL5vo7XTES8qr
Eh8nYAjbaCcnReVWo09Rd1iC8p9A+p4rSU6tNGj+MNUBmcGLA1zGDSbGO5aDmeh2QNOQT/ec5lG/
47hkdgvI1BObNyRVoPoGcWwECTosxRIpo42pQf1WUa7LAO4+oXqV1RWv8m78bmW5wpbjuOxjigqL
J7a8x49IC1fcVMd4mPOo64t7VRib3qVps/4eMeKap8OTwzRBONzIozeYpq9YA2O4oUoAoR6PoVHp
kvmmVEGM4HCsBdYhKbQgatJmyZeBZic3k0hcqVRdmGH2YiHvSFmtb3Yss2D/vAQzV5l6wxo+hcTo
yrhYvD3PpLVS1HbjpFZTYIETiRFWAw8BEmWXcsP+A1d2dND8IChlLzvnkZtmI6YyHS3M74HNP3NQ
ChMnKuxH+ngPpMy8boAglO+wU85xvgMHThwx61FrqNtnKibmMbIE1B3fyX/szF0WsQxooAjfq6dy
EAgK2EXVc7eYdTChJKZuRSdWWt0cOflIqXZ9Plh+E6DJ3RUE8jDS4XFf57GunoYe2o9FbVSpKOnB
AqL8UfjbkVmL22vQS2+bOQoCOuf0oe79fD8UZDCZLgrmD18lLP87sZdlXJekhKELWL4znuDq/dVH
z94NJyBEdOQIOfwHa7NgCaSlaV+dJtITIJ9roEzHz/AF7xm3IVW2DmG87UybrR/gRJzCxlnBbDzo
ydcOMGkQ+wiObwcziPIM+4plZaCtrgocVX5xB94n5qpMaU0rqmnTf4/74unCP7gcK0ne+bP2WlrZ
wZA/bE+NO0VuxU1RbZiHkWMqilgo26XsF7hFHAECKk17PukNEsPr5Pm7ZVNQ9drooDCSBxcCCWTT
kKUJi3ZVFfk+UkzrhEXvcdbEXV/XO8MbTsGDFUqG7ibJWokpzdkuXYVn19yITwgtk92FRaYDXYwM
GOeTjIfyMT+Jit7vCWAy9Fcpw6tZxeD5YTa6QGTh1pm46voWOYAsStxq88aSlaEDC4vueI8xAZ7S
14qDR7aU/mvOEv3CVxe8lv/ajQZ9P3OJhWurtLe0SklYiTdf4TYc+05rZZxe80MitjBtr1tBuEM3
AObaqcbTF/V3zt/IsCCrgdniJxUnVUP4EwVwa7ZSMV0AVzRAB2cThUhriQkO76svad2Dk4p/l98A
f9NhSVgBmtp0vF69x3tBQwEkbC7EO7pfZQXOK7H1z/qCFN4QIpuMtKhwId9evk6jl0VL5Vvu25O9
opuGw2JQDY0ro4cdL9GLQEOBz5DyP9HXx2EbBtzbo6LZMpcPS2lDiocWpAOv+3rbUzFfJwZJ6092
MZe9BAyvrLb8SfirM1uIdc39NTeUjaOfVN0WEg9v2r98vPPMfspJ9atL9BTTPJ1120tIn+x/6P4W
GxZL6HFm0VIxRor6dCNicpXWGJKeQ1iBQC6tWi5elTjjOinD9PgpfiPd2jWkhv9/0+4tPhDTJ6Iy
oiTdlbhNMWYvLxU8z69j7K0TXXTJZflfkErvuYSpjC3uEdjMoUqHLxUgn9Nb39rBv2MveJhnk7fK
/qheMho1+jBA781M23KR1Jjr7SfA7YPEZVP0MapEJgdxgt4zs9i3wxE8BGDupyXQO7YKDupFW+IT
RfmCGprJTDjBOBuTTPNW7TEV1se4ARo50LSfxPcw82RlI/0CAb3E5qMt9Lk9C72nLLeowqAiVYlA
ehxokdOISQCXPZ8SC1nCwaU/MAwxGYnLkQNUoeYYAl0FVA+EZcbzxVQAaIlOu0rEvCvZZLYO1jQ8
mBWu7X8FL0fZXNqUoc3trrn/VL+Xd1AlZMC3+1FplHes/lGaGdn/l+TAlEWmVqEqbw0DY29Zxj34
tsOsQ8SR5Noa37HUa9H553t5B6pzBAH+gXE1DMvoPi8egkDOguSzArMraCqa5mVwc+OMNbsQqtG4
eeyKklZ2VsbqtgIgV+MDal+LuexuGs4Up19bTsCH3TjEMAWq0HK8TWhibTdBHxF3rAeJ034gFTHc
s3f+RW3XlNk9k6hOc66+jkAykRHZ6G+hhaRAiVxdjna24WSTS+mOGuRKwZipMjwPs3AkTo7zJ5NT
VECAG8hvep1y4EqowFggNAn9zQkK4HOkrkMhsLujVx0E/X5M4kSLbI5ZU2lzXLdJwoX+ZbUyx7Bx
LejzvnkJNuQyYjXW9lwsFhGbM4xeMB9Kbswnnl3IVNESx1sdyEwouPDrpbNya4+ct0WU2T1Pi04Z
3Zjai4Kb7VJfAbEFgM75NS2yyxjdSFVsaAJiCMNS6mG2XaMprrZwfSZ+XraOG+9i28raEVqCYE3M
IoqOJu0FxmD2QFHMH5F6yBSWBQCoJftghGVCAqyEx1XIP76VktQ74jyS+kiaUWzHiuSUw7Tum+j0
NM4/UVulZ3A3xLKs64/GP7TPW+pJ/eXTA5ZGG906SrZNFhuH8UF/42D4ZRZI72LN9HmvaWn5WVQH
FOqz1S87LpDBneSjkByfJTUk3eO5Ck1SSQbKEzXwGJbdjEYdmAvnvpaVm6Roi/0Ir79ADMOmcvVC
fzH21ud8e9wOWfsSfzx+zXl3gY9p7y3Kws6xVIQIap8nFHZzuSnDB8LITF7V9KUU44ykmUltyvw0
+81vZ0co0XYHvcq1k8POaJe7oezwiy/z7jZ+CKzCB5ilfX3wdap6uCKxMFZnnk9t3iZ9DLWKdAJm
KYL9ZZF7mGNFN+2tLiJqpdljCAvMjVfzRNQoWb0bLr9NbwwuL7hJV0/BRpd28+J3UZfBHLSvlsy1
g7BDrvS1N63Eqj5VMuaV6HrS4962AjeyAh7dvg+bEtpE9o7deTpcCjhjkBRw2+By25O5T+GWwA1n
DAZvo0NRIhOD8SKQka3sX2zE5psnexL44E4p2Zhw2TMX2jSmUflI031XbY/M7q7/6bBiHSCmnlrX
rxtJ7uc5caboRoxG9vGDqUrucnsy3Y5EgiFCGLXV0lVFUmKflDuQJ2u0YgVlZStHu1a8vNfllhBq
o18EmiWrGY+jSlMwOCfZwj9TlfZZqe6a/+oYhGESWNx3FUOkFC+klSGjhDl6BNeQbya4gbF0yham
SrWWjUZsilw00GonALpyZoxeD4Nr1xb0Im4ABLySH3bJZFQRK4pia7TJ4jEihyGtb/W9BRI3CvJz
WC/9ad677nphk5WUFAVQ2Lm0TkkeC2sZbS2UYRwd9XGmmveV0aPYyDF1CBbPPoGzyoQ9wz324zAh
wXh8ok2qrMJylZAE/19YnkK95QKXKelv4wscc0gzmERoGARDODB7ucoDKv2d0PorIzfxspsV18Jz
iR5TPvIeWD28HpWeU1pQV8CJt3vjjW1b/jEaqDl7k2aOOLdM+A8+4CNxZ9uKOs/mRwxrxDog6m9o
KEv2sAKZ/SQ8KTth43fX/zbaR2rDJrtPq7IogOai2ddcOPliPDM6Dg+0bNO4BPJfLsrIDLXmCLPC
9X7lvi+FLr+51yAEGwXdrJqNVA3dxfGWT/3QUTmX6Gk3cvKwH/66LgiBiiUC57C9Xi31H6ovx7yy
eF6dGinDhhXXFSDgHD7QbRslNBVtseD6ihhuRsqqxDuaUTFj89euKz/hvXT36cQ93l2RcuCmfyBC
gzrT/6Xx1Q1867l++wzHRl5/DaiQM1Do8rvgnvhAILexbPajc2onxkRF/cpbC7vSxFncK/8l8JUm
TniiIgEKI31fft60ixjNyvAnC8ciIRvNwZEnhbg+KrENl1ZATXrHZvJeJGfnuslB/M+t9qdahkxT
jZj7fy6dswaG9wSl7V/E1NIN2Xyyus0c/mzLWZtaBYZ5wCop7248nqYZI8dfp0I5IAOpVjjIH0i4
Jnv6n550+HaNHTEf+5Gk+UDcV6leRjlfY1d9CHJ2RXfW1YkuvevdMHNCjXoLHenTV3ETQL4P79Lj
yO9CmbJTTck1qnWs2AfpvztSK2JsDaOnwt2hJjvvz7O8SN60ej59QopW1oUh6/9wmR+5aMa45qYd
fqqPkOXnXexEqPshu9a16n34CO1TgRX0zkIUEqaLAHt2SHBANff3sSPvuIugmQKiypOYJoCnA7Qw
eAyFT3iN1PDoUj0UdtDsNcFT5c18a6iGEb1YZ5ObfN4aAfJuMNV1el9UmpOODpHh1EYwZA5v9lFs
Nk5MLxLMBYWx4qH9WczoV3aE+C7EyqE8PHA7mi/Q2jAdt4ugIs/EGKOcdODciC7xyI9LlHbJGtJ+
cqsjZ9pG2NOtApiOxtJKe6Ok+WG5nKfcuiVeJysyg44R/mLi9aoyysHDeE4hSgFQrFwdDk1Pm7kH
tQ4KswabWlK+dcbD+agVhu3hfmD63ETSFdvGMeXW2+xOC/pI8aRrVN9Z1xWd263MnqQfek9qu97y
n37PApe2Jj5CDbc++kFMSRCtaeVHgpUd+y/mBHE2PHFwGsqrLMFZCLndf+xZvorr6CLtoTN8HA9p
XaDTgk1dK8zP6kSfuuTmvVt9DH7UZrDfQFPyUjpDgqohh0W7KyqKNm6wZsqs+E4cGwLe4O9mtscC
k83bUJVjD2uc4CJYCpbafqGxm0/qta6IB7pw6IaWMh52G5Q1rJSDgdju8nw3wCN2nf9gkWs9sBZ8
OW4I/HxR19cslQ9dKVV5SRFlzfteFT4rSHsChFzCQ5s5wh6tGJ0K7gbd9mqOjS3oRjaQp8C0pnUV
OIKJoAeMS0NxhLnYmy1fhIsPt/3uRCfHMk7CkKAZuYHGq4UfTTpGTjviTPmIsDOwm1sEdqiuk4K1
4Da3b9iSN3plIAn9eWENSXRIV6D62Nd9P99k08aDNxBZQT3Q8U0dLPUZh0pdkqie8y/9kWD7w4ph
p4Ca4Eo6XVqEww5sor1Jr8gRHmH/sabougGxRW+NieeMmRChFGMAfel8iWAWO1zDsrJpo/1BjY41
/VGloEkPJvZTJDBd9Ezj2FHj/D7MfX5kPLUmE/F1sWKXWg5hqNjHBqx5gxiznRfoMbgKS0Fr9PFS
+KqS3pMB/6342Ray5Y2NSYCc9BCSmkoFGJdT8HJmFly4+oNB6F2yjiZUyF7tUWqoXmihKBPA0YO8
bGm8kvNh10rZohWFIxnHkXpajb+Tw3ymnTSicPkn0UCoKuV3UYaR1t1oZwRP5qta36L8TJ/JGIbj
3htv/wfkNiVpSrPq/IyOFwZ80oYqMs89+0OJv7+n53LRxYfszKrWaIjO8xtcoFeNpOEALNI5wND6
duOUabiAQQiPoLtnk8CnYBEqLEorkFsm+irXwtCBZDde8OuBMjy6t5IkwgNTuS5uYrPI3YBb+0k1
af9rGQMUrclKRMKA/UqtkSDPQ2chZ9y6Go4HrKPoRPkJ5OCqQG6MsRKxvE6dTNWl1sp1fDcNzHeA
EooE47d1Jj9IuYr+kf5oVRG9DphGYiKxK3ehJyWfgxWTzpAXhfVTUdQJ7gzDyra8m08nqzHbiBXR
KfsVoOzZ2TDWlxUnCg7vsZd4+w1j6ZWS1ejtQoaxZp8Nv3TBurVKVVM3oJTp5IdTAdefvN2ye2ar
3pJCuO1gtxItXIl/1glbQW3xVCMN7W9EMliYOY4IzdoS42kWXMKL3+SZYfwKCvUOI0lUfL25yRsB
twi77kjmxxRhzn1BAvg9qrCDG7JG1CP3Cy6Np5ZM9T6awdjZ9LVKrJg7Y04WX2TA2UwsFQjCyBhP
XHvaCobkuVJtOzuqd4TzwfcsgTf1WHGt0kaAPWpzzD9ei+PTOsMnQ99WFujF8TtwzZH1NLaZUWZV
Ss0ZACwclcoPqnfBAqSLDY5bfnEi/BsARBAoHH5jHQNWsk4dgCSOwdMAMP00s7gfMNSjaOMtmJOl
Ggsb/RBLpCVCpGrrSpWD6xrY0v6Pnn/ajDEoPRJ8VwGAeILJdUd7NHLY33PTKWo2saHgvB0lR5cx
Q+fkQ1OfVhztUc8nkUGzlRdSGkx4fzwZyjLgxsLnV6AD8x/Z3SKjXiAZPPV9LIt3vRzxLK0JudoG
tZ+a13WllvvdUqEVyyLfkOwpgYDl0Kb4dIIXpKyP1eOPwQtskz45opVg2jMuRKRRBA7kPMixco3u
BOlElqQTkUlUahR5Gzx4T44MSEKYE6Ua3oPqJ5Web7hgs+S8gIH8Gm4UmIh+zS/kLW8GPy8gfd0/
rNQg3xYAtMR6XjnQfJxMEE9fyNzqyWbAcN/nYgwRGKHxcaGxvGNMoHK+byhBv04n/MkBym6hzZnf
JxmsM+99gANDTDiaBCvFP0q59NM5M7YHxNvvJGzzgF4C+XqyF5Otn7f+uQd8VG768JC5rSN83WME
y7jhQmbmTL9ryx41iw9g3KBDikOe95cYvRQ0WszdTmSKKFDWrhCzXF2IA1eJUw6rvLzSU8Q9cSA3
USRXr7k0bCQkOWcpMNUTYDZr68m2iC78FQcZHmhhJmVvQ2A4iT6mJD8iLz1BOVXbeD2k87LQn3Tx
3AN8ZHqqjKUuozren0cNFfunQcedaBzrabeLD9xss6X9B3T3ggQQEj92JVx/HiuetRGs6IfUlmeq
Xhao6+cHV/LpHPFfbci50oEI9bHQyMjNGg2FI63PNediFsvSQLZwPbpbloDI04wUmOvUhkhsQZP+
vX1mbiHmuPlcn4ou8kdMmgy2fnlbajGHgaE0JPq50d6Bz6VQOcIqAfrIF+XIOG1oV3xmmi69qGdX
v1AxW60XsfLUc7gf7NZkv5Dpgdpmq/gOKBNcUHR/pS/owjvmcrbg622AvKpcl0HGzdlx16ErEVaa
CdtZn6iftCDMZFuZW/VQgcu/b8BpZ3Zy/wYuVyUuP9HTf6hpg6hJGIZtqY5Dis/vlt+pNEfkgbSB
9Tpk6YF8zsAzOJs27KtVy4bolZOtLAAUp4rOJv3rW2jv54U/SkwoFq401CU/kx8JkWcNyh/kCoHw
dY1pgzBcBBgxA88+LO/khfUOjXzUOxD4Gp2cEna1wCnUPtjLoDcoOk+fjbj0mg1KoPAmKKO6nWnW
0CFLN5/XaycMNo/nVkePMGZeOcZXum2Ojcx91HOxE1zjjplbiJQmOa/qaXyXU+309J+c3g2Fq6gr
iWBPsyuaHieOpIBiOYvwYmBilRUhvvTvTv/mF7jVgA+j40z8yfcu3ZlrwKthis97u3zFKhGmMF6e
+lCUG4d80+BEK+Een1SA0Ct4070wtv44sscLYpbbSfD0ihjnb1ZYagNJyfuglHC5MgEXZ9HY/gDH
F6ffw3/B4JMuvh0pW/E3nZ9KoFSci0nC7DLgKB0siZMAd/Zo8lORjTsLHQXHfXiVFO8n+0devuMc
lcNoeqYLRrT2HOnb0lOgK5WkcTZ1FVSjqaDATMc5sB9Zo1toswCehNWTz75XPyehQD0xyhpI1JIo
7bXXm3+FmIFnZRLDVHJvPFBY2UbBvGB13F9YCOSud/urHoAMuq4Nkq+qIq6x+kk7PEsmfgZV8OJX
JUsjdsYKwpFwhRfimNM5aT2z6MKYA+RDZZfb6mTbvo0ofvMKLmiNhs8JpNbSptdkCqCdwXhe+KjI
WCFhLO3YsLlfNQkEDIvbJtACZBxVjYc92dw9ahXwxFeDkU/cFXGxMSJGUnqozVjJsnLr9Hu8H5Dz
NKgurvbtBSKU9udleMyB6o/xiBu4ZfELjEy/OeEIkOWv7167bGMb7wVoCDunEXP3RPuPUYOf8D+q
bTpj+a2SbQyvGKxym86ztrsLKXhf30pvwJa61aLEORRZ+xcgshTa+iYMDdHn3Ds862B1dQYxY4uz
EKHN4VVy/ss+7IOjvRdTl7v8ot+NLAkzMH2I3Cim0GXpE+YcnjnTdeVqKquInGOkLUu7y1gaMaBN
8tvIdIgg3ixNBXM89rDK1xjROX1qR6NBO4+utgDmV6AGWsJ6k4EQWtG9MAePE30k3taBdwjtOnHT
mbkO93PwMQSZPwDmFj+mtDIUkutC3VFe3f+OXdBD6zMHXywig/jDpAPblhSJEJYVdTSUzc/RPpg/
9D3GBN9ForN6xolc9I4aZuS/BKeaBBRSspBxA0txnygUEiM5YO1XxFRolenkcAiWDHsHgOjd06q+
A8BtZLScg5FTkY1eRZ9GkyZrnpF4u0eapN9eOFK6aeuKY9UAUyPkiKU8DjuNrpXZSJyON2s63AVN
S8CBDWpjI9HMSy8Z7CWTZibUwjHGfbR72SVUI7+P7yG6GGTFxXmsPLd74Q2TbY1sJC0GQkgNe2rA
QnipdApmOYcvMkE0OnOCYCNCqCY4lEoWK6dUC2z3cF1aouG3HjajDv2EYkI02YRvLup7ro33fH9J
XTfNkL+z8YuliSeQ92DHW+vKhf0x0klLnKRcieCJWrIp9O8trRCwD2jo2Ge7NVTGmeN0zszG08Jn
1sOkSOPuq7B2u8a91xGqOxLddVUAsn6K9O0Y2xeWmeWML1qUZCvtFR1jUMY71/QQ6Pgh79PJcFdA
w4g3hqz6rh0R6LjcaYBEq6SLWXdGlvb6rEPfyUr1xDogZYUETV6s/ACtlS9af9nwP8v7MHQB6o/5
Zsp+QFlL5E2Pg7oIdlVHm+9fgdTuPVLJwvm9mgXb2cIavk7zfTngmveFvCA17zIv2QaqpwTmKoot
Sg6aULOlkJjg5l590D3LD76mxq7uNyIwONQpFlGkv+hT1CC58PCQ5MAIq39Qq1ieFIV19rlMTzac
+8X2KjrsHev53wVL67D2g7H1mFofM6cargJC4jzngLIy7+jhfgks7zdJ7Q5HHJfZg9Qko4aBYQ9q
pc5ced20PhJH37YnfI/DiNePAou4hl1SM/x87eGjZoA2zhmr3AMezvmYn63+eGMtxVxedUdLKqKi
ciGXd2gEAVnQX2vy1woK1CsfWGWiEPUGA6Rnh2vz6brQJBmlTw83EcuYpGVMphTVBAn1PC/36ti4
JpraDVCCAH1X4Fl28M8+FXSc29VQCQe4SdFLjOyB5bObmWsaGHEgelEM9DXfdNrxDSVNHTPPyszh
RFbGX3z9zmdmoeGR5w00XBmCpHQbgmEnTAoI8PUHUpgtMV3Dqer2CdexE3kmOwYQ3l1xYd7wFENU
hHduLQO+NmV7lMXHL+3i3xueIMVncHyuiVOY8ZAU+m8v5THXz9yIamon/aAqKZGCssAoL0+EWPEg
FM9I9nYyFC5mjLRPDuz8+C4wPyxyeAXOI2mzOQrNKVjbP6B+ztWf0CHuiIEHE0u7DkBrTfYWywi/
Zd3nS0XcSOPyhKR+svA2mT5lSuOxlPquKxz2lMJ9PVcJ1ttvWrnUdB6tFIMy356VHCBxQ/3O02vq
S4NlPxq8GXMeCdOt5fZA0lynQtHhq/W/Zzc1k9lwAN+O0lvvAbcUiFK9tnebTY75DZ/vhtEMJ9jK
x5IWxZCxPDNcVhJCNXbf987E6SyGq7JneMsQXmd0DlqrqLdbZIjBxCXJ+8XjQ9Q0pr6r7uMKYw3N
WwLg/rveOTB4A+rh/j+FDX6ey4Q6TRMZJ9NrRlxdsZjfe18lA3/vYGAy5OoMstgtZpl3jxbbkAD1
XQCJJCx69rej+LtUR7ALHR68C3AmZ1turv393nXuYE9BebZ6nWDWVbEeBPWOsVKls3jQMOoduHqT
IuFSgdgubXAMsamm1qbwC31pubFH6etg+8qvJQ1CszElU9URCwORER/R121W9UTNzcU4EXvBfp0w
tJJ7ojxgrow5j6Ku8nWhBRj8DwQK3fWecd4UyBZhk49ts6/0Dg8xZ86+9pvTikn6EVGSUoc0Jfgr
vgRYHDFhqHBb/SVwdZna0rK4P+uFNYRPJG1aPYVoiaF6OzQYk7Ab5TPL6wnvaGACyi/WuNBMnlI6
AgJardVS2uxEVzAgquWlhveFEtVZGQJ3bR2ZuiNWLBdWY0eGjPp3bNKrMt83deC01cPbz7xdDPLD
bk6wSDcVL+vNEjyZ5emviEvawyio6ptmHvytvJPe6m7HAt8Ih0eX8qVuv9eYmInfkp8wArm1L8T7
6eq30OoomMlwIAWpBo50vtBNMzwRVf5lhv/WzvQV8m71LTC18x7KmAPqYenCiksgKGkeQ1GazqVp
E1z7HgDD5lbejbv5z9cGiIQHW9eZd9E/NhsUk5seQIjjvguL7fOZdeJKovLnBP+fCFt4jtLSjPAS
TuoupoZ1v73GMWmS+xeBwAy/gheEO+z9ND/CwQOx1o9eTMPdhhhmW3yKe/r41golP6oCLCfvjsIR
9j/BiBCY84q6oLK8vL02Vm5PIZi0FYgthDLM7O+gnEfQ+HP5ISh4ldplkJK3zs0X7cP3UsXkf0Bx
Tw9Dchj+kJI8HAjhtypuocS3LJHzdYW97VntQVuqrSV1/hW3FZHZgBdgzBhkS5ovEL/N3Y5rUzp7
S7BZF3wZ5ke5tXm+UiQBrw+UZUz21tIpx0ax+6ZdfN8xtsty3Y9y3NEp9IBsQhU0ItDnCWqh/7mo
DaFxwdMMj6O34b6zW5jQbb181RH8KVIJAdRvhxR3ofydlSpew1jOXOP19swLNrFTwHggwTijjq/L
lf/4u6dPTcYOZgPcuhrUslovuE78jR7jkCARjCgRntM2/CsIcTW7n/2SjBCmXCQMqbrgpt0f5Wqy
59HkaYdOJKX1hHRPYviR6t38+tc8+alXJF69RqNovJGpUsHscan9zux6xOQpWt+w/8AAxymJFXjG
ia3ssTO1avH2SyRJ0+n5zdyMAzwDXt5akETbKTv0z69cgKxK3MTNab2fkMLwYr69uvZCPh/DePaP
GjIStlVRZHmfyazeE6S7q2RhJspvRfa50Fi98ejRQsj+QzkcI56EQ64ssHokHE9fhVMsOVyqUOeK
yqVq5o4KWmLJhAZy25iBNq7Pj/X6YhBPJAN4Tw8I1NpAJGjbinc3f2jw1psTc529dtlQWKV5ZEPh
yEDxEmJpImY+z64saBQtvTk13rpFqpxveCmojKgcSB4gl666OwnUP5HwrraVNuornw2UwZ7RQCSh
sibNCwXo0zKvE1sqifDwnl8GLvMyMPt+t863xW4A2pEkJ6WpBdPxI8Wzv388eNLUJ9ZA5zOh++2d
THQ6EhpGzat0GKP4Ipdr28aWnaEP7Wx22DHO//tBj5V2Sb7LUNNkvxkq8lSu3/Lgbvp8mRMbkMfc
48lw3sGc4aI1b2F7oLVzFGLHPlwDoMR7WfVbIinTUzVfUspzatVD6YXJU520RfwbMwI7w3T2xzb7
jlTUKsM5rgtlJyBsryBsIL5sJIQMtmhyVnkHo5NtT0VgKC4svBxtJcgmBu/eZGuUGFerNSOcq9oe
BNN+Two0FMrlzEv/trK3Ky06hlKU82bV0b5n+56X7bAtr2NrfPn2DXMEbBTRr4qTETC0HK+Y3mdh
45IoLyv+5me7zOYJ2cvNHBT3ErOXQkfEorwBb6fqs+n6PsA6quUxYAj21x+J/A7fZeQroQIioJH6
GABjUOpkwPVu0ZWg92BywOyesJooxWtBmIjQE9QC23OUl0INJWzwv+XjJarlnr/LIyNsSuFgVCFQ
MJgy3CZnprdVw22szxC8rwifbVi/LchXPfc55nSjJfuJCDLFB92geWIXdEGPoIds5Xp7RNOQDPs1
aRx9906rGRvxouY3sk4nvkCZwpbyJKYw237UQFxQarjtmxTToaEMMLg5ofJOljBDkQcvdSomuBzO
52HxMud7Wce7qKwtKaOC+NMOQWuvP7Q5rqzEOE4/z1JRI8ZJyLZWwPAkBNybFJw19kkSidrgd6Gz
M5EypxPUUnZGLQKtWxjTYqoIQ2WBoM7of11onUgp7o0Y9mcMcpCbbOftn1MOnkNNAQwAYvMWaLEq
HYr2MLurlmYPKqMvuRtFkoFI5ube31qkFUgStD05MFPquIoRdIal0SMeEsORgyfAbo+ELuYASbQK
RZ9thzMglVdIzBojO8B6Jfiwmf9cFLWMtg6bRdRiYmf4jdXUbRxYF2XeDBUNhZ3s4pLqmeLjd7NX
3D8m4lxif4DGp2/uLllW1oDA8f+ObvRPmngPYAeVWe5XkO6GdGRnTJfBV7OCB4T4YWnUx5tt0FFB
fEnnqZ7n7zrjvm14l35miwGh8rfGgWb+iKj2yQHcOH71R1WnkHvdjhe8Y6R9wqDT5KzKQR2Ppe93
wngXKIpxuvdo69hkpeKI7rk9L7m+LUMVGnovBlZ1mjusT87vzvVLg3mwdmNErJgD7V370N0sOJOb
h0HsDlsrQTp82CmTzoGKlYzK/eSC7pMfqczWQ5UBY1Orx57N9eximHvOwE+pNB5uCFDCfaRZvXJe
SXRlebt26QE39P/Kd+bSZmRSt+Nw191PEzz+/A3eR1bBBHB8XV3SS82rerm2wg9KVbTZoK0EEdtC
Y2zagUcqZJGLhRtQwPFYhed5Qe/QjI/uwqW3bZmt3zL3RBjgyulldD0740RCjJImPLUDN1bh3TT1
T4wcfo/dThgmRrhCyWGoocy/MEnD2C1WHSmXd2QkPLmUSDxYgC/gGwzQDrI5OxVIDeMLE10XAaWK
6UPPsQofQLRpPwB9IHeoI9rloG8bO1Ps6ipR3fJvlzT5e3VkTeTyirxKrJKS8M052lYUfQrvbcnz
bXExiON1QjNGkfwbfDxtKc5oy8SQjru+O07oYI2nUCJfmhaS0a0Gx/z3pHhkG3ruuz7WXDVFohaM
APAxxHCNP8C+o3Dwb+1Md2a6S3BILFgCFF/EVZfqOpbrKVtWTOgoGnPJiNrx9I9a6oAuoQYyO/m/
O7Ne0tmyh88pp05gTIrZQaPGGE3p9lueE4NVAlNGvXXbei27C1QgwGmdapRdzglO0H9CXj4dGl9P
RZalBl6uZZLUzu186MYm3o0YAUbEsi3Gy+xRukQCrxCVIjb5+CEADcKOUI8sfFYtdYYbpS6khb+A
Eq0fYpDj5gnLb6V3FpgOil9KZdddjoA1NtZ7VGEevMyobL7hsUyQaOQ+Q0FxUNpc8AS8vBb+25cp
q3Ptr/AqcuIIQSu35zQyIzeKTVfs2z2WTBSJimN0f82LttrkWMExJRQKWsqaQ7uQY0Dzd/6c9Voo
Fm0GTec2Y63ihZNjer4tQAITkzLJlV7V3XQBA3Prw5v33IyEZAdralCmp0QuA7HuuZtl8aTaXijY
zzrhEYmTF3B4dcfG9+UH6oX3QLtr6E5fJBqoxROjePhKasSMEZcG+/+BeRt+cZA43TIn7iK+zwHq
1HNPudj9ywq2Scl2B0CSSVteBpMk5ejDO+19+iNB0ajhy1Dj9GsJyJMUraOSfZQWBvSybYlJ0tjq
7Udz/erRAWt6B2DUYZ1Y3OUWeEX2fGYq+Fk8SedFxMJvbENREymkYxbPOTpavVvI4vOx9dKikA3D
izLEhv5UTs5JXkPStfd/A7GhRmvZPRRw/udVAmRuFT3hf4Z2CP/7LSJCdJWXjSGEENemvPKjpAPs
CuMD7067lrJivHjcRHjbZrSUI5ElpHfaa/RmKcTYsCbaQ56SKbNPu0WSS6k1PHuOxRnZFJYeC0XK
1QDeK9bdePGfToZCFCA7/dKK+pGXMvavdCNFY/bb4atwim1sH7ZaJOAvmJZUcby+eeE6L6pAUTfS
niCL/B+KnLFKWFLuw40tkOsB45cpk1jkMa3TIjHYirx0wv/JfyAHdJ80721BsbEBrxdgNdrXIcYV
oSq+D1ThRppv1vlB8LRvm8fQyMxKcTzga3dJ1v6KK4hnTZPWEavm03lPulsrKfgEE7tVe9e9L3c6
TKPNVJoybQUVI/Zzp6YF/4kgnKv9JpL5DvJ9XYYKkrjRHODOKtxClhNs03BxhBoJhmtw8l16Ar5Y
R2kceJf3bP4TvwKKn7C89jXSldUaZ2NOLrT1ii6ZfEObde9bo2XTyoj1O6p7l80v21QNaVCoxclu
JIPWvYm+39kuGxiWbtj2ehZ5OLEp49GkiICPOkNv5k2ePZnYUoET9uf6wO3moxm5wU/evIycPOC4
5mAC0qz3E9i+p7/uRQ+iPk5j5W4eY8WvPMfTygT0NtfnULmHc3wZwhwscigKTI5mV0ArRR0hAuag
bzqvtV39opu+/IFayFxvnr5QLC20sTzivGy5ctisowuqyCet7ig1KDcBsjojdmfdWQQElRjrbP0G
ObS0PPKBnDqcH1qqszERuF2tO9Xml256npkFi2Dj1YqDo9EgPXnQHVrq2kOPj2YALDYjpRLFzixx
NoSzqcwRGwAL1K7bTLwyZEKcBJl4uI6gwu67/M6n3pWsXuBrYTZSq50jSJI5i9DVGsXGvLcBK3FT
gUzScErYrM51NQ8b0SiD8/oZJz5gVgsApc4CwMeHysm0ohIz3aYDgM/WVHzSxxTojzSL8R7AqvQs
9hSvteoGR2LnzLw1fco/5Nj91xOy9AHzwbfU1MgtseMRVJsDpWpbSlenWnr2F/085ELQ3ffRA4OB
aFORG1hCYHGZmK3eimwC1keVDgge1sNbWOSCak4tIK2y22pgzJ32dXYmv4aMFTFT0KcIWhv8/wHd
yHDCDCzw3jwS3Y0ocsgGosSrL61pOl42LOYgJOEktXjRG3br3fMHblBAfSp6Bcll9PXSWqvCczW8
HSbjPXdJgYztMS2GJ4GwBEudearOXg9K4JZ93eK/MDhEJpsZsr/DXuU6IMoOvEn3ul1aSaJ4jgGk
4HJ8zL7BEaKn6uAD/yhNaPixnj1takhLevu9sjgnDmuogScJQuDnLLRBV+af5wHiOwujp9yvk1Su
Opw1a36jmyQo5a8Cuv2+WPrc33uEiCxwMYuPXWWO1XzeSaL1Iab2cLuIRE36GdUoh/YJc3M1h2vx
xyBlLV6Lzv1E6boDspiuDYgkDB2jneXadQWRVk7aHn5eFo5/fjq/ldYS46YV5UoDlod3uDrbARWw
2r2eMDNn32hn41bkTAJXGKD1oqBwdF1fstZy69J7fbMyybEJwoJB/07QZTShAFU7r9WaSX1THIyu
XkKi/y7LeBlsXKk7EDJnIVjyxmz3dehb7c82Zr2lLEA2wYftOT6kZ8mP6I+7HOGiNPs5zGXDGS8s
l+OS6OkiWuqApxTaTL2PCP2RbbFGb2+4E6CBNOQp6UR9PpTos61WLt3omigqK3phV+M3qtRegQBN
hpSZBgEeGBChnpmxsbcmJjEN7yhUHJLV4vQ+PGqG37RsqB3XAwBsZ4Imo31UxfW5AzGgz948g+CI
N4TJMmucTiUrbV1UoHJH8qoN+2cFnei3B6Jk5s0nT08EK7cnhpQyZymWQGFs7kTVBVuvyF7LPGT/
Y4hbef/kToqT9O1HM3A48JF3KRkOG9pRjT1chJBC7yOkS9PyvrI/psEcxi3FiIdgcIADnoncY8Sh
ilzPLQc7d/+xYolV4q1EY6Jz0rCVw2WTW88UDZKkKimuVm2R/YJrd7BnU+j/4CenYNRTf8n5avTC
zVwar8L8M4e1eh0S/vObDooc3gthIYi3ujnL3/hagIFBhI2QEgDpgG7TUDWw7waElVN8oKaqJSeQ
xeJ1ZGYE5foxyUo9nJNHUkJATe43Iw07CGw1s/L6bbzGA6ix1yD/UMLkmbxs3iCc5g/+exzMvCHF
gj1rMVxT+X0FidAiR9eZn4benA4WbPPVtF6xWS1lRO0iIc9mqMnClGQSwaxWppGzfJUCl94h3BI5
oLUt6S/WcY1qttS2dje5mm0taQpYlMF5lJBQAOG3J1/X4POvP17DVHiXrlh9V/S8XKsSbS4tgtHi
Bi+UlJ7KKntJUJ2ZouIDamjZTmCGPfFy1qsukBCovsCx+CRF5tHfhcRILgWu9W4NsyE9KwcHLd3n
lbI1YTJqcConxzwzxTACBC1dVB1Gra4CnP5S3AFvuGBOHBXvZFejekd3OnQE2Tbsgx9ycG+1NV3g
pveVaFOxTYoGPJh9Tyd0MymwgLgeqsMEcrnG6/IkQv2tMEvh4BKseapjmmvLGhdCeZH+czuIZbeQ
epOxIMBvE8KenCXwUFRxgDEhA1WYiQ87qz6Trukz5G0A/JrCn7aQ3j4oSIoV9cDCvsq3ZgUwTioh
tMsUvQmdmjI0C8LGbwVwguGYaEuPP1y5q7vRXYodTh1492qYEkjW7rbuz4k1M4U+Z5Tw5REV/e0Q
fo6TRNVwQUNN24w7QQW/q6PAuyTjCwW2vo1AhbPloXXMc+XOTMBtSuoQSCsZCuXpazuqDkxu3MfA
dtrrILRF2JvcgxA3rP0LYMuAGxyRlivfMRqEeJUtt+3nNc9J3HKo+YW8/OKwCBtCkGV442kOmOk+
8+O0MJQPFrztS2Ffjr4Doz5eh14YMBjqhRS0poMUpn/ftFlTbShrnmbe4QXvAjnz1Xs69gwMx195
QZ88LlB6kIHKRp3p/v/JLrv0MI94h9JItwZ34dWXnmDGwj7BsCWkEJ2o4CdELIAPmZOc86vG1I75
Pp/CGCIgvaTlqorE7Hlmns3Oj0xukbuPc1tmWhKU8LZ+rdGFAl6Do0bTybNr6AzufXRmswgyTKP9
lBcw7IkO6KT6WhbSWbQZf4QHa+dJpQVblPG/zMTWirCtHxf6SXk0B4yeFgzFs2YlUjm8VV20CPCT
UfobhzFHHMr7PkdIypYRqmyq9OOv4svMQQatNP1zoHPMY3Sx1ienrYrID+fPtPTxK2AZL/SzV2l+
xXxWG4XLUlArfpQYjSiO0hJQsL1k3rWOxu4rXV5Z0M6VHsuv2/oUkuN9B37to3GkEwIb5E9ZNgYO
v0C8bV/4nxBotBx+r3d9aUiP4rhNyWeI4dDO/VqF83dd4aKVkVT0RBEOkyKHKgR+YO/BqsJ6ETBc
7YZq9DmO3KmT1AWRO9PlFs8X+zFHEZQvV5oTDZQGBAu+QJ0UYp7YRUvQ5NIL9C4YBRxfbDNW5oOj
pp25TaqcIgY9BV5L2RyLl28+u1nqj/oY01ioCFAShUHrQM7toIcuicF3oNCLMJhMWQvZ9U8Q36AG
+BPjJlQlK8mMBQ6D4Cfq7S8G00Ags/yXi2jwj4FRVLYdywTRzq7rR5xn9piQ+eCnaGiSGkzNDJGw
+10DV+/8hYVfSIQYrVSszb72OAVbqP/8H4zGZOXziXgIdSRS7HG1AVOD45LJP9lq095MuJkhfbi6
164ai4O58GALCJbRmv34TUiLNmz451JWRXEfEXMXRWum5sLkYsAEuN5zfmAb5QqSZRWN35bEKTEo
Xbgh8/UtDVQdLATUEyN4FwAGx1hMihIpX5p/dePKparkyp090MXTbyKWDqjXdDsjF/1CMmlOHi9J
ZPDwiLpEFIULdbPzSaV2j+JItJ/l+0fZl2lhCHQ4AENAeieDy+FXm4Mvr+NK71ziNRgMz/IUl+6f
WncHY971LW8IkCt/yDf4iUt1UfcVTkDWitCYcDdRQ+r7rfR+0sJtoLftfTySqFwcT2iN6iRJRuS3
zFdMp3RRahDArovMquNF7Psu/Db6X1RgzoHVl8HbGofRS9lvflTr0nXbRHJc7mdfxv1ERlvAvIEA
gFyipLRX3bhwBBfy+T0XQ5chROtf4uRIHjl/Eh4wYHweBjUFcD+jYUMCe5ji91WM4l/6QfV+vR4H
oyO0Tvb/WaMA1qT/UBb+aMwc/Sq9dKfd0aGL+DAqYlGSXxvC2GWZBnY8m2PUIIJSxxXa6ok67TmR
Y5UL/UdseNyFgkB2G+UdDR1PSylO5Y4hO+hukJR/ngrcQh+eX8rj7T/ab2gEM7DQw1yq0hyJcyyx
0eenu4AhgdTANrisT4D1Hp4n8W7nirkowtkcWVJu/se+YLWeiJMB5CGkf6bk+i7x8gFV+uNbT/aW
FTVzI859EXzQIfE4/bfxxNmesgnZqHUYdA9dau/8TaaSFcEm4kuEUdTdLvJp+LkZDvCLb5A9DLCw
FXMxVRhL2S8ZMp7omQdeJDekF5zu5ncBWRzhtQvmzUf7BrLDcryEW6fEAhzqOssCca4yZYbG02yZ
OSyoj5y75mHpgodA7dkUBR2mA1AnRh6qBjxBdR8cNNT9uVuvKyTN2dPyJe4LDkopzIq3jI/j2SH/
HWwK66anbFPXo5kppMENBc2iO57QmZlYfi/sBwIDDewquakuRqg07olJK/tGwURdBxGmPHd27bvn
hqKt6rmdNzLQ1kCj/bu36eU0UQxEdCieRekhAyPMWeVcgTffAjM4y7Wud4imfZU+XXem3iS7ShTf
OEjTQGsAVwCWiDkqVIllJiCtgbJAc6cmgB+jT3+LATd7Klt/9efgRFmDCRo7Zb7GnpaHbgZ8HGRH
ArQ8l9CgWX/BczblvEnIx0pl2Rj4tPtCNEobPkF8N9wuRlKhA98lyD/wyfEVYOSu3oKSFXOs3hAq
dPEbWTDXLruEFKtTwvhQB863e0egBTSDmMKRZSsC0CNY4HioFyG/+O2P3bAv47JCSD84cUD02fBB
mh9ifB8TxBM6n21Q1zdlgTDUa0DDFk18gU5rdMPE/Iq0AGIdSs2mJjopWiyVBr7b/f8ogSxdWKIW
LrJeBPlB8Dg646vusYkbOaT7S3ivv+QMHmnyiC7CmRw2s9acRpgzT8yafwmKx2IqEMXILPSMagXu
vCYb+VxTpRZnuRrjHqlQERMe1marL/BszbLe1CQYxBvwM9eiMd/MGclGzV6Du7dITvrmIt4Jx1/e
DGYW0fZZHInixjes1HsbOdKSfYBfV9e8ShHTMxcjaeVQ8BZdfcHgeap8ul1v47kOEhpDin4zD6p+
ge6GuY+TzzkcQWxlT9f/H02oFRKLHxuymqhSNRvMtGh3UvP0p7n603TdFm84LWSgjNTfS79bLRLp
oAnXlQycuO650gvCLsDxyoZDirSRJMxn5k8p27Gvim4QVIVKmDLEc6ZnJKniYJ4BKcUi5Ew8i4a5
82jDB+qcR3CkOfzD1YfD8COTSBZI8pLLGZfqxO5ySyOH85yttQ+ztSEBrw+PVcxkzhQlhz1bzc8v
f7Nn+xaw1ziUxW42Z86LecTsDtrH4y6m1D4IzH7ch7LkYXjxL9OHz7A5IcnHNdBsUZWXDO7U2aIl
WGXYwVu4/ZGM2qPxC/s7M24qM5Bw2/dK7Rc2UfgxEsNBqRZ40rIojjZOPRRPqxsXw+DDEvPAHkMf
58SHkKFmZcEzoisO9v9fUzvhUkdFY1Fx+3sMCwmJJvPTz4SyjW2V5F+TN110RLs+Ch+ZgmO2irNi
rMOCXNWL4nSlVSCkMieKN4/EXkkKGVhImBxWs2s4UHiPBS6HExG4r0xEBCX/fPymGR7POYIE1Ajb
8wQIkqpRTu4cU32is5bkIZPZLcRy3wufriqIJKtZgUImMOP5+ro0LuPY9NN8wPXrYTZ/5FheMwrb
n6F9fw5bc7wR62MyQ04RviPOXGwqQrAxKpv6sfUmpeuVEXLGSNg4WnNCD8nxBeoAPLI2Qqsgs9Bc
ZiTJfNqlBnoizD5bHb6x+AozkC2A9fUdpLA4UbjDzY2PAKENkMMHaPvTr9doX0uhfPgLO/8xF5mX
3LLRMKYBt6PTBQ5ezMwHEmF1QVPEYSUzYXC78nwfSpOwBPPi09cpEcsrXdNtifRkJ/GGGn6ligqJ
pMrgFfrPtaQYjt7ZaadRbP/2ramqZhhkZiSKMz0uu5GJAa4Rx7PnrUcuJPZ7E68RoH+VBZkKsaHg
ulRcVlOS9c9oNg5G8MAxqaoGuLmqb275ImAwyxu1K8md5HIOcYp0BiNGM3WVOs07qpV3yZuY6MzZ
8VfqcrkSjIFbXsZNWI8kEmRvquBgBQ23w8A0ZYfv14P8qoZEOku+114ZTVpfdxrmoE4x3UI8oszX
btN0Hraem5kgrutKk9apuHc2uQtz1k5dVCR57yoTCelXo/U4Ago3Wg8RMh5b4LUm9zmMSl9D3Uq6
gGeKSX8p8SKajGAUGtq1HCK7nMnOc5vTEuJ+ZyRhyYclXxYqHl58hJ1HwLRbY2GEWrswTBHmrAf3
XzeGD1oz6ikzzotb8fPiLp7Fk8jWbq6redh9hLVFjvM4Z63d5qB56KQdsNfsBmkorHibPEeVxPzY
BoHZe/8SYeFqBW5+j3o3CqZixUXTCCFFmLSg3+b85IybVlHlnIS8vtBxt4pXJHC9m4mTe9/4obBH
/P7gZZNMIvviGptfxUrsTxgqHTyEypa8GKDHtiRARqG5PuoXTWZYa1y51iEOUknlZXiY2oMsVfk2
1+eWZnq1lq6l4hZNIXeIVFmTh/wJoDQE0+5j6sMtWtC3zkk3BKH/GPGESMnnueGCyAwexAZXi2lQ
0aJxIjzv2O7DheTrVNN6PsbsHiOecmDgR5ifjeZQ38YSjRSmt0Vbhq64B4QtnrN8HTWv2UFjBFYb
wvwJVj4Ql/jqH59+GvbIzvUxoSVKKGzNcvniAIkpGdXW1MDVc9qjmxWmGTPU1tjKTF3Yf45OsZhs
X8xVNldS+wLtGVFBuTTIcsuMLH8tc8w1d0dGIjBe308j03iXCbXKSC+cTAtT+b/UdBx7JViDg57g
klB/bcaMThj1TuxMgME71MoljDhj8ALbpBof+AA1IaqpbiljysKWjgHVaBwhqP2UBPdVRgG2yweW
SbqEhXMSGZdRhjGtxyEpybopuM3Bz3JLgSSi0aLj9Dj1xAUpxojGFBFhibnI7iLIxIa9qXrrQAKK
e7LWLzaQ+Z1iByKRoLH5WvJQpcAg53lcHvQpdQsgKPEPBJRVW2Vny98b40TEtvROIACdZHZ/hifm
gKbK3egUeqQLY1X7JPJ+vHOZMj7lp1yZzGQIkh0RzOf/YKRVEKFt78aRMP+TeWDNuvA4OcDlXB3g
7RcP9m7aaMnGT8Ck6g/7ZooXeoxZugp2nU99bu073c+4/RiGfpIhgrWNGvK2b9dFYGEZ8IsM0qm6
6MsjkGgrU+T5A/yrV2CplZXC8n0V76JO27Y2mTjQh2TYClvGFP2+EWW3xIBxjSMZOSW+6FtYdLgr
CAikIw3O7EB5EHcpgeTTiX+j/ZzwNdWNpK6Ans+773RBcy1AMfHCIBWEM0x6F9WyxaMw4Wsj4lUx
9qL5jhF5/BQvRAyZ0DViYafn49vf1OiNOVdUCW1YRYN/qIVdNHNxlTp+Mxnug52eYtwFYTYQgNqX
a1aNF+KRMRUaq/zMCpbX3T/gzz5QWbRtjPFzTv9eV7XUggUE/u4UwwNTuocblJFDqLtjmB2bSZmi
R0yW0EQRj9o/Oy1upwI61FehoYYcK7Mc0YBpjYGS55w1dRNKA0yf2oWLEYlXJOLeGgzwKDoP347N
2akPmfHcGPiUnQ9Ut3hJI6A2DGZ5j5xcYud90CqmmJYivSjeuDDfvay3ELqMRkQR3wMPMCjTz46X
6xA+RhIFhWFT2jyLR99hgxe+/WogU7q6tWEDO/CitANvgpXXnZ3C/8VGalQCzysZv+rOw+1FckHj
9PZdyJMq70dqQo4oBGTyWl0rnw+g5xljMvmf7RWexUekkTSJEBJi12VxxFxJLtvwYskTmtDUkgCk
vhc/nQikzQvNrTyvxsI9GpQccIlpTMqhux/u39hByhYE9SNVUvTA1ZLKHFfWpfVrKO0IWOjm+0rm
M68xqXUvQEaswdmGpniCpyxQkpVGLA6RWEQ9lT4mC2zgaivfpwz6VYUZHJ1H1ChZwiE5h8J6Jmln
rBpJiSYgxb0DEDXlWtOpO7o8u9+r1fuqh615aWx8Wy9VvQUT0yy+rRc/uoUuQcfKReDi3K9Q7bwW
CcWGjMs8/uMWOotRFDwPLpGfP0GxNIcFsDDUBXcBwMMgMV7i+Zc258E0/GkuDoqxxsbmO3Ph0jFZ
pMVV/rGdbmhXfj/7h2mAggJdphP1Q8S90XWLgeovfrLZ8Glt98QgHrS/tOYQ0jVLchKpw70OU+eM
ly3s8Ungxl4S0jyNX7oSbCzjiEzLoTDEhFVvglbNmEwIc8PBi2RQfREPKKO6AQNIAYtKh4QPMAfv
dHJ6hJb8WBSvu/pTYn1J3IinyUYvARB9P3CEoOg+106BirhXZTJRbS/QtSX5KEMz5/HmZf/s7RrC
JI65obbWMLI2fhR7FJJAmCiW9E8MdJnAyP1NeZRBw8ErgdxgRE3KBk3bzqzyanVu78m2u6x3Wr4D
ZSorZ2jQ2rfmtI2pNN8LlmVmXVt8M9/lOJuGbrhxbTmAAQkwPtitAxgmX4YnHqQtDfg1d+5ULY8j
KKs5BaKyBvNGYFP86XQX95QAHUST10p1NTub5whWn5YVQwLzj+NpelXvCG/EChrvlvFZirvPRf7W
xsm9X1AK9Sj+h2GgGjUARN/lgb5veNIRmg2saMNSYYyihoUTMlD8sPiNch+y0pmk4ee/rtkqXFRl
B1ZAWG3khTA/NDvzmYwaioBtKkWmMLT1FuwUQMDNOdJg9AOedVhv0GRvyoih6k0HtEj58C0Md+dm
72uR9wZQoHMSm8owtkATnvTjEOYgLA/HegqowBL9CeK0tuA+Yo3d/10hfR00UB7ipPEAh4PdpQfu
LU3zqa7i+qxdeMRfaps1sjB9OpadA365hveI9ZXotEpIN2t9N4tD6wmTuN/q4BIm15D4hRLAxRRM
2NgK700EDyy2PNK7x5sx6tapJm0R+fz7xKu1dv66dSABU5R3bXx10h14BW94/wK7aUo7qxKskphk
luu1M+ZygApViYrbCLMMKOFqHmjUu0aOmJ6XYZmr1gEoIW5neuxjEKk5TODkDtvGZiDuTmjYuT2T
PeDVjUyLf6Yk3Nu605NuVcva0aZKfyzUxlSZp0feytRuB1yJ8O/5xz/p8rR3qvU9F+yV/wYwCSfb
4Zg25KNEbA39bqecCrEy5BDyIcGeH0HknIDDsLVEKA3t5tJMlVhXjRgIOyvDsJ5wQ95hMW7lnYUJ
CNx4O5RTMQovGMi1WlS/easXYgeXjAyVidT7wlMu76RRCh4qEhQpxxhAtRuQHZl2WzO3UeNU3zxh
aRTsL5oqibuLnGNRQLIgFj6i0sqRTHVLROq5r7UR44S5DLTEwlEtFAcPlVxYL8NPMIRMlrqiBNq1
DOfZfeB1udHu5Wkusci5Ew0uaW9BuuqAfpTDIEVGsbBQn9ecln7fkf6IrwKCYhJ8+nt3M2rVkfd8
zsgnmNgVt4KIkRMo6anMCNRkblKbWLg/5G0Glo69Eoql1fP6B9qOW9UPWDSrI9jApq4rTNictoJX
thg00LdjsfZpxoxDuBp9Ls5ToIsgd47DXx/3qmjTNkF3yNinBYYGTWjIIyYdWyu/ZwONV47a2QQ+
kqVKS8b5Ccw5lcDo53eMZgxu4canzbZ2cg7I3kyGvmqlQ/XKGllWfeO42nkAOHVYcLv/OAlXFv05
KlvXjtqKBV5Kxuu0TfTImHAY9VbVLKIjYTNm01iz40GGBlx+N24eGCQmv/DrA0hhrh6/fVhhuqm4
7x1s1WyaVumGYLXs1DGaXsvW7zqjeZPmwxX9igmQH2RE6VVL7L//thUMLMBS7SNqPkCsHLCSApjZ
MGcTCmr9JbI5X3T2zRprjYPjEg7ydN0Dj1AweH1unnymaT4CymXAS60vIpqRSWAi4dwfdkCN66i5
aWmrEg8VfA38y9l5B4w5hnjVqTQMaD0+OJUhaWDZ3GA3zxecq23jzVRuBi5xqB25a47eBMG9NmKC
zw6pI/jU5VCMOM8OjR4b0eZm8f5WMf2B6f2lIxn9bAzMDrutn7jjOuq9hTYJplE+FjEv+r/7sJmi
7hw2O9yYTK4S5Fl5/XcQP7ZD8qmArHV1YVAcVuHl7uQrM69VMp7rqN4Xntk9crxQDK47G4Ijq8+k
LRAPJa++kByh19dXh2tMd0JdmHxwCNPa78RzNkzhJbmImGiwpwU8O3wPf+4RG6MoJV3EvAU4J1a5
zHz68NRyIX0vfRwU0I41mZoMAjTmdFnr12zrFMRnCXVSQDeiQhhXZ44vTAANz/952aonavoQ1zzR
RTGhOyvWCLj93KVpo4K4YQaRxgag8phtSWB2vXJs24BVMtP8qRTNCSmkCNE0flE0SeH2tByxw4E/
CrKzE1UqyyQsBvQPDUJelOXlKVfcTW3lBpFLRKMUgsb0KxxBU9IwCbSjnlqpj9p8gR4NbQFJHUGr
YRX+BVG13wo/ym/5Y9RSorOo+NvKzMIr4ifJ1+At3xd6XMTIFoZTaFG4sIbOaNLImsnzyg5KHH6K
wzl75jDdYP1s4s25oZAx9JquUqoWqC6cIMw9KIlGogYb3O9I5ihFJkUYnsgEAJAtWNmEMTmYLMbz
xEkOngw0TbZKuskY63HitN5SbEJUzuLYX+B9NLCrnlYjs4Mt4o9yc9DYyLR5mmtWv+mIGxBHPqmr
H9r2txlRRWVNQPQZB75jzGhTDdLLN2oOoc0s2ElGURUNLun2Rk82fbp9tZ4nVX3pF0Ut3BHdof5z
fylw/+Fq7v3oQoN1nlwzVi0q7yMUVTjyakL48kr5GwyrUYIKTUEZAsjgR10gcvXXW0zNCD+X+p/7
mGjoQ4Zq9fo2uE5JgFs/VhZL6/UF/rh+xrntfeuRPChwV2zV/pzDA45/v5pvhGFOxU+gSXj4E23C
Cky2m7SWaYbiWx6o4y1Jk8RV9tEgpWL3vw9F0oPDELSa9lZEMlBqrr7vqvuNl5M7Ak9tv5YEFMQ8
0DH0Agcfk4AWdNcuB6tFP3c1RHIfRBYfj1UzVIIpFYWD7FIJNazjct+G12SIDPWVUPg5WQJfG6pF
Jr/rx1yaCQOVcuEJp9LBqgwTG67lOLU6PcJiNAHVa1/DrtmxSTc4Fri12Qj8GYtXJ3Ao+acxD9nt
aWaKiEfQ3b3mDyxefvrf0LP96k2dR/cA9G+fMIEju9jiMgKMaBNtFQ3NOeWonmn9NXQR0B4OnzWd
CimbitjdBzGBWgpql+lnwqDOOKN9Oo2a+7jxNPXt2q+UhsdY4FcOA7dUBelet7DUHdDhzrwphUuF
pr/HrhSsoa0E2LzS81uKP0HW2aipvaaBE1rXcFciapfxR1H+Vjt4uraurvVIelMEUaztkmKVLO8z
fzt4vDIGj7vKa9hgUUxlI0q6lEBBAXejbIk8fNQW9cB/EC/LPgk/r6ZC3rGoSBnxvRGyAuexD9Lv
tlbEHiNRKosK4+St2QGO3MAnfFntTzpQCodDXg0fIQC0JVuhy3qLLP4q9sZeItKBVxowZ+HyQWE0
YCHYVA4NAo5ogFqhrY7esDaZKlsaSgvdHqZOPHQNtBCGRZOBIQb3yoqiuxuwem2zKFcqDJGbksTE
xdY8RRh+iapezwn5oa3/bfA6NnXJoDi6yIKQuw+CBFCHQNaDI371EHMSFW8XI2Yw1UNnkQ1UKsqF
mFsDd5DuCEvga2O7V9IMQE8cxPk4D+qpGL8NgWpXFoawk0v3N3XRjTwjx4ARlfwRp7Jno8AJPj1j
MywcBV+KxloBaDuX27neiSKRCLqTd6299V/3JUp+4LSUARxO2cAWYXHS2OEDSx4yZzZUr9ekRgOf
M7iNHEzY01lgbZWX5zO1cJP+DPKfoZerXbkJbUuxXet9A+CmMEWmbfAZA8B+HDz8hxdqYdmpIhyf
hMN2FJ36KrfYuL9/2kJCWjb+OHZfXWt08PdQvizOVpzt0QcDWjFEpCZmuLBQUSWfo57/atSP9Q2r
54PYj/4hE2UUBznFLst3gxDFaTTQKYpICV360uYAF3QUAMln4A5ZS/bPfU8KCSGJaACaRzrOGBLk
gcBjT4UUuxGw5HLEQLOEr1QKIxGrnAa/iBqhxruXKWVtwm7naHQDv9jK6TXl067UFNqXDibd20sM
94F1x64eEAwGcp9HIhpYeUoJNDFVyBggpC5sZIbD7wpnlfVC3My8WldeUG1npIqz6+SbGbsxvb2F
P4zy2ziYRSCAfo089QFKrz8AnLAOBejcnTJXt+TLTo3brZlrKmX2GFnhtu5SaqtV5g74uh4ilf+6
53Cn4sMisgkR/F+4MgMrou5oeYpplrzACGUybAcCbAh9PKc2ZCOWef/r4I8QhvUMgw2/+h3lgt1J
U8XaXdA8gB6PXT1L8YbwA9e/lWjAiYtZjI2Delp3CTK1CRmtJGHhiLxY8vp+tmNP0cHh2OQ0Q64n
Vn2Dve6GVOrtO8kwAaMBf9niPn2zstgj5QEYaZ5eSVna0dZveLTRT7N+G/P+dOjHjJ/FYD4UrKYb
Nu9A3dA+HhPlmAduYBggFQIgL5Ucssv0GaTPG5u5+OxchCS/Vmz3NQfvwCafFy42qmIPqOAcunq5
3uhQN6EjARL1h7tWmjDvBJWq+Il8BbI3HTHIrc7NVnk4B6PSncVykzBevKEcS/oGASnzbg5nRj1F
ai+bajE8Cw/kjZC2/MG5QFYxxsaQ6f2nasYNDPcy+VefAaS9ht6Fj14rGkeD68rDY6Fvpamq8Y+E
0MhLZz6TFDH6aRGPNzzyP2gnItHRkczzEjGM5Y8VJbFS9Gn0B0rgBcCISLmBT/ygHqgzdya+6Qs6
VMHUp1WpTGHNr6fKI0flfX2/5VBbiYpyEGCVpneGplaLMbtTBxzcN6cs1TDIHbl8veU/6b6GJ+Db
/eQmDzCECnhtX/tstc9QL+25/RCXHue2e/IyFL0B6nr9OweQOHfS3DRxzPPIB+AINjNQgD1A0rpd
g81HrngawxuwYe4wZDiaHrvuhi7o4ZUPBRSSc8VmYNvjHazlAj8t4VawnbkbQAjO/+oD67AskUht
fvd6ylNb/YSKgrRYcvEwaWlCiazmI0+jYPcV0BKhUoyb009UdzEMbQkXVXybkJYL9xIC6dEM9Rw5
4EnRIh/ivUz3L1IhtqLI4PEoFniUwOp7fhAuTqC3hIXnbz6rsis0rZ5kQRZ1XtjVRlymQIaII0Ux
yOgvpwAJR0ClSo1DGGvMn2aXoBTYAm8FAeKpDyjkZrxbhN0yroS0EE/ee1EHGDC8T2sMF49IL0Oi
nUdOq8Ab7SJJoVuK/v1FdSuIghaR8w92l19bjEd8rMzn/UoweisQZpbBGl4vxJu58DYxc/5SAm/e
l3F3h1gcTaAFwYD97QvZRAg52zjoOKyK8ZB/ZTfuuBSLRxwrLbPbnOV/J6TAN13PmqgCd7kCZiQR
8OAfqCWVgCOmWhXGD/Oe7r50zCV8ep4cLJw9uKsvzwMRHSJumf48/igELYtllJ9dGM/Qa1hyQrJ/
PUgkBxGXWafLw7nWiak2ciU01xbsmuZw0r31mcQF5shlUYbCoXwU/BlieORa8AROakGxJWp0OvjT
ycfS+KPlwdmHWtt4kuHPDYZHpBZ/NqYzkrILmwGUzyNEIVO/l4TTWolT0h2GzTtNJnlv8DpptChH
DvgRiRHo5yUB6WQUI0+DEdmNEJYRWEm6bG73UOHMuzPpqZ23RBfnRHIS5RztyC+RdVTEeOpx/xcE
9RItVTZ4iYVZgV+CPhOOIgL7bcGCyQT7gK1F5OaBIJopVPk710gFkPiRZI1awJwMJOnCQFdebV8+
UbwvW8wgpQD333cPN+fBiz/6RrZ1I4sMC6mZ+44tVH/OIehj3eMiLrtZeddQzw+jdMCoYeMxqyNd
dwOfUG2fYLXdBpAQq3Eyt60MKTyI5iDOipXJPaqWq6wchV3DQcf/3LjlfY/OeoymDY9FTAJl885r
CCbDLNYaf8oUwR/yEFNyatPBV9stqbCYJwTmK/fEMhkrwxqRA3K3Q3Fp6KcXB17eskt2S6LXQAYO
EYWdQqixQQGIARnaHZDawXDjXp7TfEHndtn330gWLqMGuQ+puQM9jhYF5Njo0NbOmAenCPbQFWIW
xHOkt3u1hfWQLY66A5Ij25tFG83waLgiwGUJfU2c45p70QG8Ol7dzg9+EOu4bQ0JyPzS/1UHlJba
U166TTTLUe8ZIPTj3dOg7AXncCXaEVs/28Lf048+jwm7neA7zc9YSOq9in3Il8vPnUhjlqxKlKk8
cf40HInQmNY/i1WOaU7gQNFJfFsAMjIxX5RAC5boZz8Tw8+uBJDFMN3LQFNXFXXZau4HhN/0mboX
if1ceXofRLRKSlSfBwIOHdWbNe38AFKlBVrlaiFfVL0TkCD3jwfOR9pjrwentYYygKyLGpEuc6wj
Rw1ZmMA2oKPqlBN69VKPwjI4kKn7lKzcZ7TR3Os/eeMV4boWiAHqqeAQji8NKrVuiYgCO0+b9SKB
r4dAxQXeF7aLy3+GIYUQRT/iYyKk0PrkpXe9pWM/cX+X2JHGuNXUXP0VrmA43NF40vm2gWaZQL4s
gr+jRaB+FWJke9vgpNIGl4m1LyNpdK5YrwCa9d9Ts2+3iFyMb6LIt2dGmnXBY70AwuRczUm1ploP
85/SDYLLRaKHouj+87pWAi4cSX4HYUIs+EzseeoAedtujHDBo/Mbg0fvMbCIIVPjWbkOPoAM3UYT
/kXSSG1tZTHpd94HAw0wudxK2625TQ2O4/3rv5xrF6oaGzI7eXr1pKy7LvBlEsNqp3PT9mHf7uWj
Jj/bfTybZovvgKgMXtnRRcg7rxN3E+8xYO475wwCxxEWlpgkURtlQIvagknZo8SUoGwq/Wf5Kk4a
Q+if38GnJggkctrTI0u35fucu1j7keZpYOOPYm4OhIBaOHOiimPg/TIbdPFtZZZUW/dWRCqfHPdJ
VWQHXxdvkyAWBImjGQJsvqPkVf88iQB6Xi3qsYsDcc/TQBUXVVIVDRP2cRkY+O/QweaDcJ6ps1Mi
MtPX1jj2ZVYBkmlWrHGPr6DKQruy4+20OFd1DB/auFcM8UPBKFaiF40qUJ3HUnIhfOiv8iSK0bKl
hz0b26IrLDOzjDM4Levvuj37zByUw9wROXe3+aKqPFWEyU8K/c12hcQTnSg0FY83BeOmIvwxSNAg
+iL6BeHNo56YPpIyOZB5FN9/TjXhSBp6F40yg+O3OfMF6Em8+lawh/B0pfrZIREQOLYBERoDMZHH
OwBOjCc+zzzf0geyhWbWVyWKhen8kFNljNo9HZd+OiDQV+qmqKFm/hrLM5m8voSNaww5qb+ICewA
rO2Ql2fOpJ8LV2Z7fsrvlUqjuZKujhfh09/zYqzxbIbsANaJrnvtCgEqgwxy5Cf9b3Wq1qs2ruLm
R/aurdaSCXv8bZaZTd/Pxg/dUR9lNDahbjDmxE15dvPXBYIQLYTIrRAuB8UU+u9hRicJLL95q19Q
Zj1ncphzu5H9Rvn79Kdg8pvIY477pcfCctLYSVyWfVGc3J5bkKqfEyTkmKGd6IOdFl1FsuFiDi8Y
c6EXyVxO/U3p29iwIakbjM632Plo6Ca6/RTL4Gz7MUIZnE+0IGfzU5wZmuZnXsU2a7IIpLdCi9QZ
nOMksjpR0l/xt3IMF1uPmKpeEzw/nHMVX66PT02OnE9jxU66fSv9nciQ0zKeTBOW++t1rjCy7QA3
JGyWbq3Dk5qFYY0Xa5ioODVs3fyNNDV8QV5vhVxn7Rg4MxwJaZp7296shVYOulmhxXl+PCKrEgHn
LEDEzGuQuZQYhCwnCvAD4CKJyU1lO7V9J4LA3VnvWBfzMCzxp6qFAwRMPav2Z4LpWK4Cu9m1aR2e
SqW8Su/wSAsauqpnSKeMcrNRDmtC1oMdXt4VbhFNBz3ZaDO2xNVKCvTLK/gsLe5L1isT2QZVIRm7
KYxFQRMS1hLuR5Y75s6rTfcB1t97lfJLdO4vVYHAnN8IP59JIXqSjSjUb9Ymb3/k1wuoCLsjhJGp
kJjCHeP83oBFBvYts1EZRNot0lCprhtabtAGNkuw1d3InrGu1x04MJsAZa1D7jQwO38hx15632Wl
vXBZNIX8kZNsQBN8Hi+jULBoSV+05gftOrm7UR11MaeX42erl5J3k84EJ/ZDD6BrdcqpEwm8zJKI
8Y/vMllICgsGsdzg/mJy1YaLCn6ErcziqXB2vmUnghFMePTo/H4x6Gxrfho428O/phehTzgHH/rh
voE8maEWLun4/6EWuyQrpritggCm1oD6QSw/DmGYYIa6jvpeQ+14qtK0gtHQer3mQ6v8UJtBA/xm
eQHD4lrYYkYRE0RQ7MLXw3dRZp/8aeyEaZ6eyYzgDnbw5ehiIMShoOgpcx0rTzBJWSwZ01Rv8Vuz
LodBnKAcRYGKxQeHY9ReqhkXjwhfKuNCtYxIcepomCKNjx4zgmva5RTGXAqquklVpRYHpeUlNmCP
QPGYTnz+lPFs6ZvW/CmASCabuXsJYz1w5/B6jCodOsgTOT1n4iCQAjKpJPF3sHsyxYLL6HxsM0Ao
9ZCVVL17PFpm00AkZKMnXlQytc0gwJWniuz9bHHpLQtG5Vs5YBRzrxOmgJ/XeD0K6RWu5bKEYZZ0
sA3w5yUvgQbjjPq6J/3AiF1e+9xbk4g8XevQ8qT8xhYOkhrRXAGYntRyhIvEYMT8gWw2JYDaAFVV
5jF5jVTLS8/uPGCnPzRitKGh4KI+LnfMLr9XiMknpQ2sZV3sty0yJMkw+0X3Y56P/6iV4srA5yxx
xIWV2BFNzlaf6VmJCLsQEUKSMv7wfy5wPXYkFUs7nCSmRb15PKds1Pq7Rws2mw58Dx+uw/so3zFU
YjOjQ8wrH2P2m1ZJvE887HCkvx6SL99qGIkyguReKmYUw7iyMr1rc9PmQB5yq2ALvt1T/CdhGLUK
qM2chV+/gsICx5D4C4G/ditDpVvXAHwI1utXqiK69qiwm7j+1xnuesTTHzbZpvEAiFZGvIDVKUJW
6v4T0m2EarcWoT5omSmtuV8fFgSIh4FVMYOasiDDr9+kZW05N7t9c9oP4N4i2XiZ6z0lAZcn584l
L4SBqvD7f1I9EUqHEOcD3ZGPFMxZqe7UoB3e8XG3KTmZC2QdftB8WKoKmYBxcQYmm284CBKIOtXz
XXcZfF25bI8RrUKSGVkTlm15Ua8XzDHSAzYAcWvm4DZIAFVkgaVAXPD8BuG7jvPCbLt4kE99OT7Y
6ivRimgYJ+b44ur6lPXK2FM14Od9GEritQ0wXLqWYCFHXpiULoNGU/etGPfHbXIBNGDPmqWNlZqO
2D6lxn/LnTBN1NST2qN1R7twDv37xTBiD9+xICVpp2HiZvbfLmP8ReiioAuSXnlrJYY/IzJC7D3+
Wjb7P9/bMWpNvy52rhwb6CZLLhoyvMk3wUs/pMSDnn4gC7dbIX2t6Aq0QDOAZTiBBQJGqilD/zJG
4ZvuniuO7bnQI09fxltQKM5xyGr67EW0LtWyA1ChYiF547OsyOjjeBx4CyTN8vbV9IV5taLutZSk
TopPCFWxB4641nGLe7SMuK6jVahiEZPLpGJjmbd5fcJ+0hNc23qISmEmRaz2Z3H94IzJH+i/4HiJ
GuD1qB4z1JPt7LUAPKTDX7YDqZMySo49wIjW93zQ1/W464G1e/2RbGpSQtTyvN4TUauH14V1wEdc
ZQijDaAsZ3wLYdftHwPtGGdmLnYEEHpuyP8wLQ7b+jFXOdSHiadCNIGFsJdRgOgsv2kHbowvmMQS
G+WykW7mF7XhNOvHuHycC0tilg8XOwE+vUEd6/ofYWa5qyfhlWZUFB1/st16SevuFZUeMLxfvbd0
JA4vv95wkU6xFX6BqbXFO+QYZGIQ3rYB6nWiVGqV8QhbN31mKDN23is24moy/AnthikUFQxQTGhY
6cEDvc9MbzOLieBJ871+NyVKHFsnfYVjcbD/4SNX92NQ4B6x4kJz4SZx/7w3x7vtQs5DynP/9D1+
7S8EQq2sHU3/GxtG3/Bm6EJIV3cMgwrfv8Y8bfNt4vwrBRK/umxtJ/pz2efeFDIdEIlhdjwRDbZO
s8RMj1ZAPTrTZDA3bFz2Fk3CXRS7tzgNghAe4uuOLgCRfc9xSRWwgrrzcA2Aw1GAnPhoSapg0u0+
l7HU2ZN19TqqVEeOT2uIvEFV81nEGX2PalcPi6rgCjsBF2LrEpIAio5oQ6O4fXAZYCB3uYDYPUYx
YISUdNL0axpzlbewud/iIcT7rb4Pe1Z8vyW+721OWNZ/I4IrdLY+vseSvAmFlUNDUkRlLhCSIibb
ujVZdStMp2O3ST46IW6eW8kbNX7HHV3J5UZyMFEkhtGOcMRlrnW2pN+52pO9PCHE4JiC2FEE+5cx
gJXwoJv7qKJS83ptE3iBa27eUstRab/+qQvXM+lSAXEkRsKT0CVzjgK1w5rQF7E6eM8wIQeqFjci
rwmsXsI/tVMiuDvzg0GYXqPPGHH1I5KJnjJBluvx1O0C0cSogJetQ2LJ5Wi3rUpo5rv5bg4hwjez
9vYb96g3LxqPenAmB2zrIs4o2FrdR4+QH5YQuunSrAt4agvhPWgCBY1SwSKMWZ/sFJVXlsX7USeM
P7z6rDcsbCFjKn/QCiHR54arW4+AzQ6SjPBogj6Il3QmcJuP3kfbxGfv67aa3tGoDtaIvgKvqDY0
DwtkdzwkL3PgEzq9WN5lwCyY4EveWsjXUpCSgXB1UMBjRwrYRkvgHx5OhF1Ros9PLQ0HO4NydSjq
09SR1+BFGQOyxeygImGH+6jc11a1d+DB60iJKB6MHr/aMn3I+yOJLhQ+Dng+4NkIcH8pccSHNtbH
Ss81ZPCMxe0KZtOG22epDuWM5n6o8aGjJGMg3PN/JVKnKR8Zkj9xC17UupajxHRuOJfDmB8Ta4Ny
8WJ9P0BDHPWTiMjdjHQ5NLxsU4SjD0jENDeaD+eRj1bS0wJ708VHLj2CDOt3u92c4iCBftKXd0g6
pqyz0u5irFMG6+soMwO62Qqz3Y17iu/83GWSNMcU2wFnbOVIHIPUbJt4W+UQuO9B0HebWy3IHOSX
w5OasmBX5FnKGmz5J3w+bZWi12Yf8iv8yYNYH9WwrhQalyiju45MMdpYLBXtSOCz2wUlb5q+S1TI
DNgWrh32zJVnvVlyE5nVNZMNpByOCJPuUbDsTDKIN4WkuXADiz52Kw+sZUYUIBNzU85SizN7YbOg
EbsXXMlgdP33kVP8vzid+CWd/a1y/MlV8AvNQNBlWpSYrQx/BozRB+imY9cnP0iDU0ZpfwiUODQv
DusRds2d/G/93sU6O5Ifcsni8wrTL1OeudPXuWLhWJd55MQhfSziP5tpKv7SWtvR61xqWlQwnZc3
UOM6Ns1qKtOoGhF/WemEA3RahopC7YmWnPvgkOLhjxFlakJzT6dixigXracWYCjdDN0Ls1wzPMBK
6Cxs4TAo4Fh2AlOVDJSuNE9EN77FwmseNMnNdAzcx6xGocysgeGvlfAkEUl/IAxodo7ojZYuiKyG
BZwCXJLyZp1om3PtZzMyGKVAUr7Uqgwx1S6djbUzr/TBHroybQRyMAbnE6GOtszzvxFTzz5xr2Nk
aHmgp12ykhGFBFGp00xAispU20sOVd8Xe/C7mqQ83vmKG2x9Yz2rHH+goqQ3McvOlpR+R7c1yGtG
nMGkJv7BhxXXGPJjngnhe6QG0VCuZntt+m2h/GmzRJJ79wBmAWbKoVTfsgQFvzbWgnHgao6ZYwp6
ZTnpdBB7nSE6u691dD15/AEvUHgAfSRTVZZfF/bL8jl0+VzMXlo9BBVklarzzg2XWA3vWGpk33qX
LuyPAg20Ngzy+M4H0WV8wOP5JMohcQlvLSgaPUpGl+3pXqsFTkljgfT1QK0S7Zj2ACEs2vuldMyQ
mWlHAIe5YXGnLT0ftNNJSAI6NDrZlRTWWBmdQFOEFPQax53UkkYxbXXl5RSD+L3V2mmzTYczQ2C0
S1BvXPXJdNcDx0gWsApcsVDKe8rEzoIGy5jfeorpH2B7VBILGR0LXvQYOJzHiT13R7L5qm9w4yh0
UpcdUdw5BalkdIoIpS0k9TIGQHaxNRmBuCnRTb7o9A69Jccar0KblYwGdnQ6Oqc+3JiC/KK8X6M8
tZmFJFEB6EyGixICKJxxBIEDcZpBJYFRDtMCNsNc5HKi6OZ6Fy0kfEz7s9Sp1weatoCoD/pNs98x
j58RHGYwoBsriozk89dT9NSFHNoSI+blNhn5Thug7777sw+ocwCr1PYOpOMVfCztowA+zKZVg0du
5HA4PoBrKY2bht/j7JmSle7RU+2LkPec2zzH7RZtbXBv5foh770CoGbwZ5oh1oUGCaWEj/auA4to
5vFFDTyHWB6V95ofsJIM//4/12/40+lPH2eYqjyy+0U7RURNB0cs3xHffaMuZ2cyuKQUJ7SPmAyr
IOsjDfPEodYO+6Fl2IovFWEau0Prf0mJUro17YP89CxSCjgMsE2tf8YOmfQmPEoKZNy4G6aeU4U2
nz5KFeWmNpX4AQ7nviI7pXMVboRk1EnFjjmWNhXQsWT5IcewCNjqvA6zZdxv3GMOrU4viPUwPbZ5
vA/BrZjsZL1BiMqY3KdxBN0P9QTvlz4bNBMS/2Ai5Bt6uoc0jCHtFLs/H6j25W4nvb1eJKEDTSUY
Nl+ZLmFjvC0U6dE/RuzyjZzetkTNw0O/eI5H1Xi/7dJ14FAkbsPwZvzb1iRhEjw7rJpN+V9G5QiE
ajv9kxQvPNmL2rFOtvhZlszuBUIiuZu7rnpR+rljQO/GOF/CUrJuMcgNaul0qbRgjU9lxXxIwOED
DoCyB2nmVplKQS7v/6zkodebLW3pOhMnmJm19neUThrxelzTxrUhsmxeOESKeOOhSmW+mvpcgYn0
1YX3ECigi7zLjAqW/yg0eoVHEHKETuwoLGQsFsZPsDE8SfWnFKkVhNR9HYF21aopCz32//ininJU
EZJ/TPOx4PE+xl+n6dvTqIbwF5TbzaOfntg8fPDgZzDeSfOhrwxGCGvKiuZAEZW26KPdfnPPd5XK
JU9Hi7Y057dn4MWiZdpVX65/wTITBV7AyuNQwaXkkD7SLQTKoVmbFnB9Wtf34ISqPppEibtjfnSo
fVtDRmWsVaa0fe3qTBRNgTYCYaGqvxhCZ3w6hD/tslftY5Md0M3w3rxeAjNksgyVbTQ010x8yqv3
G1HeaGtbm4akupYW2dh1qXek11LPnSnVkgMhA5pNCzOLyoVxUdydUS4ZPvLv5YgaWMiAM7dEYhJk
uyzq5c/WEnfzllABS6CvR/PlEOPuNMJqczbJzo0UWjXh+YTtuKBUnw3KBXXydh0Ci4g5rRuUF78Y
0c+GIq2sul2TzXvlAWeqi3e3YDV9ob5cfr58Pq5BY9J5lk6iS1SaplRXXfTRsUiHrZgM6aYCnZG1
kM0GBoBNT9gbzY0swLyC8OkL6rZM3QEXXIjJlOb74VM5kwuaI35oEmozBELmYNtT3JCGkidRaq3P
YeraG2p+fCIBzogaYw/ZIhigIOWi/chlXCk45U2k4PGulFMRDg6qnVtikyps2k2Vue4hxdIfOsYv
cL1Fa+0XchxFReMq0CgiOMalbTnk/wKTJ/3QCbM9MpSYDDvfMcmKuafZulfo6qRO/y36Kot7xiv0
cOqrSoHzHXZeT90W+lnTUquJsKWNMRDXGGBhSWdxvj0X9BigtPABC+axYRQo31z9bGEfqIOraFiA
Cr799E4P4Vo36ByKEC0IL6LqiDWEXqRJ/tJp1qXwGLxwV+0xqVirKwC9Tl0EqOgr/mdTcol5vhvD
ABUV5ErP3ycQUUtqERYCqxuq6dF6C1M/9CxV0AFOtYNZfdnDEJcl102ITFoGlVMULVqx9DJwXYtL
53W2gWO24mvq1Hu7BiAvTjltkyrHocKVtKp+GTQN7z+22yMlnOf+4iqxzeQmUOFmINZr6KsjGqdS
QnURJ4kb1xxWDyF7zV7q+N2dqldyadJcwWKDRnkovIKh7RlrPHKVz/akhIMoDNUOfTxdKcC4S76h
F8l7OsWKxatH0N3+lRD7uxOzCq4DN2il96ZvoaOLcvoYaqbiQyyyWpdrRApAQv/TgPSMPj0kBVOF
Q3YPKG2/AQz+Vkh3fR4/HKDBmnKInRdkUZfVdSQGqEs9Ppy/THwqW0i41qpIMYguUoenx9zNR0BU
g/rzR8g8h29hLFt4xqpZLjs/5BQkLgCYONzzKk5TanZvAIAmmefqTFJAfIyhIRps+qmzUMFjnuj0
mRvOQcvrqDPnl8XWuRmJXYTN0xSw7va8aiUK5Hxdmqhrc9l7/kFAZewzWkFFpTrjZ69zCJKYmNC8
2liduVi5B/WdS0r0hQ2vuXk3DdASdAbuoZx9Hq2yAa039Bpb4gJuZ19QK77N3XH1B1cIT1HEnJss
9tXgFq3r9qVT40qz6TKPP+OdnqXnQP8qPa5meyu9+TowAS6kQsKy7uCDaIg008juNpkZnthpgdRw
IhIPl7XifjT5rRIFV8/IVnCvSJhFi8fzeTTWpSAeoI0BEAT2lpwhDgVeXkOpzC0wv6DZnClkLHBN
nkqEHNHpsjpMRqqFRNFWjzREXyGKmJFDr2KEf1U5VwJJvsvNdJB84H4twJqZhjffkEDMj7Yl6Drz
SvSEWhp6F04DFM8vGTMExTTrEs1/w95AQYd9e7fwXrG5svT35RIAYwhb6QACYmro6b1qmOTLMHZl
+lYzNRRTrtTsMaL/K+j6b7NtioSKCPhrZk8FyrRjTFdlVWtxEeqvvUVM3qYON2ZZSIe7irpIUq0k
pKdu3NeKt258eU71CQC3CdaPMJXNPN2Cz5L8GBZjzpV5O002/iJCA7OKzWDHAfWZD2IFzbIMqhOz
v4uQWuc9mjCQnBu6sc2Ubke67REdoJq74ju+GnMLqjrLtVXU2EqUydmwIdZ0/rU+E3k76LmI+RTk
66GwpdVS0GBhl9pmcgYoQMDe/PpBp9CqTVCeh1ht5YSQjxRrHpUTS8cRKiVDKABiVdTwLmddK7zj
LcW3C0cmYVPyXiaxoeEtmwzX7Tz6hcPEHoL/wn25TxeGNWoKZZjChv3YmVskCaRm+3CGoUX9zEgm
KB8S490Y9Gm/7DrFsluqdOzHxd1csKqnXp1GLAqO0iMUygdnGn8zl6TGSrv4OccOL8NbJPPJFSRd
1x0DaSosAZgfRj1JdHkPstmzxrz6Ac1cfEPDUobp3i/cicuOCl4dXZpqPUoNiVKmQsXQhmp9ABKr
x5pcINVDNQrX4QJ+hQVKY+YmgiBim0H0eyxYQRQFI1p3m5dJpSj3EdsgYhUxwRVlFfAnspdxgdtq
S5WE4KY52DpkUiBBzfMsSEiJHg7JJnvHAW1bZuTd1KWaCwnAznPdaWP6PQ0h75W0TCuDR4yFmDBg
JkhGm2y6K0SITz+A3s1CDukNuKmpXdQo678bxovu7TL2Duip6BGAO6PxT81a5E6hE4kdq6bhfJwH
N3/l2qNWnHmY+Gzks0Pv/W9F/+ijdM8eWuEBsIOsQOMC21QWhAOlCvFSb4aybQLzydQy7n923upP
VY7dY1OCqtI016oErbyRVZVHhEiARbEzOT2ZdhtezNyB4hmuOGhV0hVUMFtZEwkVjIwVsNokMOfD
M0IpB9DfAT9OfzJXqyD/44ovXLxP537GqhbgX+h+0etcrmRRXRP5heRMDIpCfIEDcp/FjYsHiTtE
oQu0HouPFkEsO15Z5y35ql0nmO8nD/9cCRihtEj6Vf7deCGOlgxR7OTUyyMYl+6j64m0lgZBlI5E
dqCdPHS5Sw6UZ2NsdlbndRN1rg5Kq4iuuC0PMLF6X40cVrgEwymicGp3bHKG+n5nrdrqJgDmxRBI
k6qi9NbWUL2nrn7W/LOg77C/2ePyHAwpj84Qt2DQkp365ui7oy7umuBKYDqrt0ycl6kAiwUWAGuW
VE9LNv/e2xKtvX2NQoVX5/RhoNbf07YK9GtKI2MuIFAl7PxKCrME0Ew+SUPtRChqXYi2gQ91BeSl
ZynvqFjiLE+1IOkUjQBcfWip4dYjjSLCrdFHX/+UOO30UKttNJDRIzuD1fctfjdKynnbwMvtWWeg
+brp5an8NipbaJFGVFbIwIBDTgI8l6cD6e2nK2h4H6XaT9boXtu8lZf8wTD9M4Y98sCkMY/q0T9e
aQYiupvIo0BuPQA321i1TarDrmOk9j9b7e7PXMCQbDJWkL8Xwo2uzUXCcKmrbU2yCtjCcS73j+3B
qp4v9JVYgu+k9R3uMPTOcWXkcdKke+vSZABzH04AEyRAyDjBgm1AOkh+I4I81cZKo/I4KzxpDSdB
o/jOVQbtwBBZW7MZeHbiuXoVGO4xisBRnp7doQo0P72UwtE/x2Y67vcWeEFA1sX83qyB9JFFf7u1
N17RkPK/Z/Hd2i+4id278/0JgaI2GSnxMLUpf0fhmDGIbdq2WR3eCkAGhcynMz0UjffIsJusKIKm
UcycyWXjjECgua0nwKQ+k/mMtkSnn0rEbuXNVKiy6OG8fE8SLvA31NQZtNdN3OLoX0/idixlWs/4
NT1NWL303mDTRduUearJk2nZioQFT2YfwobZVEUVLp19h6XcUuSS3GOjcR8l3X9WI+mpPRxrNdg9
RrkMWAl+V3BHS3g9ZHxkpTsh4FrhQuae+3xwSz453avU3g+yS5xeTO0ZNR6C8n/nPfRZA8RVyNuh
4YcWRqLO/b5TmAQ5lpGJjcWgR4w+KupYnKKa1M6+si6HXh53U/yWsqBn2CP6gZig3keRnvdkRlla
5hszDrP21PjZIARTylIRQXAO3oxywZTaYBG6bB0wdIuP/fEgrB4fDckIXmHECqzRE3b2J3vB7NQt
bKO5781WYWEOgbWxvlocl5TzEA68DZPnzJYHcTjmjC+QocMhB4zA3xyMfPpENBj/2kOjTdGQ8fSQ
9Ko5bcLv2gyns1QYe5vih1YF7/s930uYZAQp9oVTsoE6X7xMqgb4vWzlVSUMKjgnsYZ3/jnipDRB
FSpdYtdSs4MEafzInbpd1RN4uP+U/fNe9yCy2l8X7z0YYXS3mpRU4MZ7LAOREJC2eepWs4cvsTw9
/bCsNpA9jvN0o/ypHcTSnfdnsZf7oa9AvSUvOhgwC/x6ze9dRgh8xDZgSrpO711TsI4a4IwCvFqb
l3P1G/np9Yrqx0a70xf4d/tVhiGEHlgpORHPnIpuGppukwbgBKc914DkuoyXAJXNWF2PpoiUJRZz
Os/SKJiuZb1YQ7YrJo6tUwczh+Fmx1cp3yHR4JxsjUix/t1tHPUXAWk565R+ZGa2BzFcj8oT+TxI
KNs8NvI66Eh7YGuflVrfijAwPjGsbNfsvkFJY3ajSMBqTf/UO/2qJ5KF9HykkDMdp2agAkF6TTAz
+hBm/1jf6jOnXxPu4tzvu6l6Ng18LGCKzFosi+wCUBnSY4bncukwoa/gNjcuvc4Mp+BBbD6DF+K8
ogoCqAfFKoKoZ7gRUuF9YYx7GKGQOuJd7bWLxkD03NK/pJCjuPrsjvNGnHOi0r8brVIlZPQWSNKD
SaknR87NyX04CDwY4qHbHuKn4oOA5m1dWJnGpjQ43Fm5ymNNIfxQbGqfl+JS7Zydnfl+dqjlVPXi
/cNxZ/8BpWeQ/xeA/AQqiBUoGSODR7CwOeUQgIn+HmhiNMe2NEfdmWtcNMo3HzE2fdBckN4npyLV
cuJRIPafx+QfBw2wAN/MAQW9LFn2g3JW/aHUwbrA1+hG5C0ZHch1QvknBL3nFFcX+sEs9+QJnVnM
UYVEmR7wszKrZB8oA20o2K82MffopTLKGt9XbMwI2Co55Zudc8Q2DipyYqOgleYbX4Rm8yt6CDp6
CMRvSk2RWOHJlLeCrr/lhyb3fC0giVyP7EDFlW4pICLTpN8nriy3kNbLJWW6V/lfjgFyJ9jGI2eZ
16O1sIzuWGnSdfKBCmkFLjXPSK3USM6fHSGlA4YZzyqqYtu32UqT3WOl2Xy+v+16760AUUpCtET4
V5lhEHzApMMoA3nOlhXMxX0j8xNtgpZmJ9XjRPXnstAhbZh8erLb1uTkW2O/NLlk76qn4WyDSJwd
bZ3DVRLvyk52yrQUwUwmCLx0nJI2nEexdFroVoqD3cvP+LL9t5S50sut83ZrUWBWJ0Fu4XlXsS5l
IV2pCTUX8NvHE0UaNNxvzexuNvjU5Yh3oyJoNaMJ74KGzFCS3SPgMUO98NJS21kpBzlVNbjncx5/
rOuDI2efv5dX9NnzCjdStJGpib9+AgOpekvbsdBG+JogKepdvovAahb3Gm6/cAEBpQhHNIBAlpEl
w0Kmw4UyC2WSwa/o8rD8uuNS+pSOD4mFTX28Dh9pi8L+X9fcNPdHPFNnW1F9Wc7j4qdU0xotI4QE
5muCi/YXwlPGP9fGZvd7bhl5QFSBpyjlafs3A65wus2N9mV7mK0cq3lOmy922sgbj3THsHqP3yN2
x3wmU0I8ZShJcKbDPq8/SKfCabNx1+gfrZt60vMu1dOzJXTY/lZ40wa2tAkzxBYbAKHEfoxTsQRk
vglNmXtS/HJZw9RE+Ol8hDKXlBj9psGnmbWjawryfTZfisjOndI+lW7hB1kF9AOO6nTdbv1NwYMW
AHMkBk08AmVS+iZCeaQqxqjpLCQWLSlFzDzPE8p4+hrSNwRTqFBpFfLSqQKthEEDcdE1JX7ybLNr
3P0R2l7rxTCWQwqJpD8vz08hcxn/Rrt685kUjLF8SE1YOxul8T/VWbu7IwyDUtct4oTBb1wUMcZd
vrEDDZxjuXUpb6alRohIdAOw3R4bV+Vc9SgnI88yO9TkDD/ACO9lnq3QWHI1SY5Zxv0RBO4LBNLm
B9+OWFBw/tlFBNBNrOnI9viu8oopbOP0GGY/ktT+5cg3vJeHXpyWq3FtiS29NqLVjwlOjKjWYMV1
W4Pv8MbQNlHKKsSw1fR1NiqnS/JCeK5D+XLeE4eE7llnqtQNPyQx/piIW+htHIie6g6QhLhYRxib
Ejo3kauHD2gToiylzTkCEGXYbNU2Towwo7LQ7y3x5LVH0cYqE2vpHSTpzwnaqGflLXJfWvmYoFC2
MZEv8svuTg/dVIn6z2yxBJab4D+DQYj9hCxfbPAxw7J85AGM7dlsxzMUmSGYxpTMkMLZsWR+jSvN
QtP8InkWEsShQx7rve3hBOLfRQa6OGk/RUuCx3V54xwyUOQOQlIgXV1niz9dQAHC2RCneG3u/jp+
ibcNi3TF4SY7CGLWsMEIUA20ijdCdLIfenJiislXR+r7r2iGB3Hr6UuIeMfKF8HGETS7pIJumdSG
xkuL1qh6ookn6dzXlcyLJMA79WZdmp674+pJBJqlVKyzO1pp9d9m65CIl1l3oq8StryJTZlwZ5Ah
KSem9KB+ewlNXYPisZiuD82cl9b9eoB8g9JubmTo0i3O2Uy/0WwKVKMwEsAFPndb+VzzVHwwxIFH
wvdTJEmtwA0gdPVaFI09FzS47GpKUFj11891vQazSZkrMU+6A7qCXQ0QWLINXomax+TYT6C5ANRU
8qwCnB+FITO/dXbwcyYj9hNL+MGbXP74XiiNIsZ9fhzfH7npq/bEI4714mOpM4wBZiwWzB7poTxP
Yf5m8rDWCaXPEq3DkFepUDUqNUj06iWiXM8PNsXJVhTkPL57CG18dp8kQeo6AqZ9isV1LZG0GQ20
qdilKLEgmuUk3GaT2yB3cFIBO2cZoyapi5hGNO8rgnyI522LuhTS01tCrrz9CHcmtu9x8+Gk1leg
UgkE8keaUsGI9vKPw/ev/rWfcqCAmDqi9U2fDele7xZoZ0QxcFmSmOYs2CevOl0LA1UoCsNckJvl
9bKOAmkJGffpux5N9MAKXDBvsX4mSJKmbrjxGRhNhIBsX0C7IqFG31xGV0DqDdh5aQdN2K/6XOEz
z7wvbKqEkH/ITp7uoWDJeeQaD5D917VM0R6dBuY65q6QsS5+e8DruVDgB7jDzxnmBT3iqEEbcOc0
7mXbw9XkKWjaHkzMsGzcQh50IXh6RYb99Uwx18OW9ROX9e92TPuTUlHhZXsts1vqQQ0chJt+Yh+h
ZEfZLg9aNCy/O8mZPZFSgTcqOkkP4XN1AbhOJaRBuDsxzdiSAikQ1G8Ehyf4I9See1m/J+7HlDrT
oYashfi5DhINH5IyMtLp/guSWmrPHu1RAzpIhXnWVRCDIMZlF1rwm/3xPwAdniUODltZieIfJ7KZ
J2rzJlhT8u+juNoOF0PSj2/mESfnM8SWuzFf7CMrFnrkhmyDPYGARVKrAy91BuwMk4wUoxZcwHBu
MPj5ctWrY0j6yVU9DP8kkibDu3DkxrdzM78/lEUgXetcVf7UZJPCfXAY30wM4vm56GYrmFsx7m8M
NysqvjzUxXIjRFOiyor8VmeSOy05fcVVmO309AU36aoi8evQUV4NJGOwmEDRj2MyYVBZxtYrszNt
X6Mc7tqFq4q2ad5X2ZVw/p1fA0tkOoR/nO1V7dNxUVxzE85lywSdCH8i570Bjdw1XzGK9QX3osAs
3MskpWXRGTHIL+kmx8d2e15N9MZ5dFMoPGioklJf74z93F1RkgMcJzOl4xdCsrvi6iUnEPwRAob9
eTljuPzpu+EByz4QGADEjRRUSBwdtIZMSn50WJiRrFzC+Lk2AbjGkOmUdiImAxarE8kuftkpHbFq
n+n9rgKAu4PV40NIhdfBDyEf0k3Jze3cpUXCLbJ0C9sfTEOBpFxDjtm2/bEUM0kg1ufQLILPtJ8e
AjJQ3DUtz+nhZdqk9NRsFWY0aIKhpo3Z9cBIeld3MTMjNUBJqlMA/pUtodP79RAwYhrA9DZYCsNk
d8OIy1ztMlOP/RFruxKfJITKiVvnC1+sADXWjf5A9z1gP/A9BH5qPdzHEkNpT4CC9L2Ito+faQZ6
llsTs5yKp7/MheOU0MgM9QgxbBUNWa/d/ss19f49nWW7Kt/SVlkLx2xVa7CknDTHrZK30qBG+L8B
3K4ibJlzNh+FovQ65fEYq/1bfyQcXQLRrv/2O8Lu2XDo0xxlNZKvl8gJaGOJimj0cQ8hFg8dkUqR
0nxy08zwjF6HtPmJgqnTo92bpGsBYzlxD184nPNNoaBcoML47D4+V9PMhwwNoxCqUWw6J19wEqIR
Fmh1AuikN5mXOBcTG6rZw+z0LlLFnUaW8+B9c/DyFT5UCJI672jEkMgZB0ugogbdBsH0W1OzwLhr
XGb+42a4jA9iT33oCXF2pRVfIzNWwSEJ48YTtExVPnzb0tvrqlgZFJ5s4zSYVK+TawDwJVRNZ8hl
n4zfR9/IOhM0QSsvZmGhTGGLVhaRjtviIxKaMJ8SHsNtCDQFT+l8DixmB327xCiAFV2xybBGeVXg
3HLDzWqFIySwq+rnSTwLjw+L0Dk4v+UtFi6Da/YZhrQSfOqMHSnZRQLCQgWxbKbpPfx/PwHH28An
bYchGcN8s354hERz0casr1nkzOwyXA7v6me3A6SoQFhZ1yXlwAUPC5zcvSHPjs9y8K1JlC80bxdP
j7XWgEp07ufK3NPsn1za1+zveebSwVDbkKJ85fl59+/1B7o35ijebaL2d2mBEivPBbBGYDXntvHd
X+/XuuR3OeN76O3CfHaz2G6kCe8Fy8NRAtFbaFwQUKLclSVt+JrS+hkxTAoIvprlxpwaCBOCnwpI
VIB2mS+yf+xqgiSG/ZvMdwtZRCDzoMi+Dhpc2t7z03+Qy+Yin6pJ20AKiXpqvAJhLpOD9UppZ9ml
Zw5DMWow1OxKOfCsxgDexKW9kFiYBXhWHeNcCS5aN0cOMOdejaAn7Xx1yc6H346YFKIPsquiBl2S
CvgBJ796NjFq1A/qtSE4wmtG1OBBY7nVuzL3saRsjPDdbHGMrn9J2enH1IFVLpZXbRHsAFpeQqZA
bZ6SOpZj1XxG0AmN95OaJ5Hh3MiBqLrRd8QBRVsGfXZAS+UExvkH/QDkteJ75LJ/AtQhsPOxskju
LAz7ixEtFsvlfUFbWkhfzdwbZa/3XI4Ow577j43228O1P2cZjZh0/Bmkt7cofgJkS/NnbgS90OzB
05RtOnkUGtY4kFjr4EwJTkNYycAviLIq4cOIdBydz7MtLy47mmA8DhE20dQAOKsCTU4GwLHQlaQZ
ImlaMvKQ5YLxjg7qPFWkUmibsIrcRlQ2k3hiT044nmYPPMZoW+r3CVHbBAp3QXEoiIZnzKRSau0q
cdhlJ51uhJ1l65cNLQrKzCxawnz2UltkpF9MwyqVY4DbWJrDgHFTsS301i+iSaobbkN5U2YmfQiC
gY++UuIwCzoi4uXz6/8N37Xtb78bverN+rFAWbHbQSt7ynSG0mMA7AqxseyzaO/FG2tOihLqAAKd
etWwcOZrMvoGyBlNfRJSLGhPaWT0SkdHcrOi+lRH9CbXbrE2oQd7hKCW4P32ouAbg/ec7g95+FoF
E25YQFCac7jfRMOAvcLwJKA3S+BnSWBYplh7jUEp++V03aKvDIIQL1SAqYy/5QSM/alDzXpEwpjE
OZGNWcoFc0Mz0bRmKb32AuSAHT7AhE3ln3+sFrf++pA55CiNKbd5vMnEgVQKYRefkeKWWmB5JFvI
fT471Eudu0pzgXgZlQdL+EUk/1ThWv4VNplZD/QvQ31ooZ6E9phze4qI89r0YG+LuYLzYVoQFVqW
8mq6g2Ysrk1qIALT2p+7QX4HVUaLFmG70iIhqBftKnpMahRlaih25sI2Q7ocdzZGY+zEWcwvo3lD
CMadn5T4M1E6rnjGnAzd5S/NAX9CBdJl0zaFGDIC5tusmZ6SYSUz2eyRsrYoE4lTpYcqz9J7qxVi
8tXSAHUpG8DiAsl835n9uMzCLOlpTGeqaVauu8n1qyUwmnHc0CBQx+pvVnm6qLTrcwyH1qLjSr5D
yDSCofyU767v6cQFHm1nYEVM6H6a68OxgUxCiCOsI9t4phBR+j8b8WVYxDhdNthvB2QI+s3TKOdk
r825TDOLfeIuya4S+5g0NIsmORAz8R9i6fmSnEcjgOUPm9aWNQ4EwpvXbaCF5uEOfglf4G85WHMC
giRnXSHEr7oNhZ38tJ1993/6I6J8FkMkpE4JWi7ioVwCA4zgNfNwZm9etIH7dDEHgG7w0xnTd1H8
J7RC0tQObiG9k6KcJtPZqHEcU1eQUuQvomx2OvZPcxdL+f3zDVlHHebvSOT0NVfKJ+I5U6gobBbp
m6I8UGBTqZ47LoK7pojCFGS4TlxC4ryO3EAC6xi2GNcydG54sGmt6EouoJuqoMFCRhZz+1/xsoIX
01UAZ64/Y+LPfBnBOL5OOADXGZj0zaUzGYgZBJ6NFu1XJ429Dcy/GAyJCFEQS1ixCWQDrGCVhYZf
Tt8oh257efwwU3jTviLozPhQUGra9vi+i4RSQqRFq2Gq4oou7AKRxSD9cXQYuTuBxbUQhCMnUQ2Y
l5Ov+pH7VSnjJrM94CWPc7WuOjoDfc5ryID48x/X5yjZsn2Id3UWRuCWg5QiUbNS6+t632zQnvjm
xfP/spD7hBDEK2FGl8c/41WioyFnArUWwbhJ0AEVJnzwrlaY46Ql78KiRAo3rv3J8A7W5EMTNV52
ltrbWTl+V0EyL6iqho+K3uMviwVB4U/rqEbsYE65G5rNwn/OqFMVoRYiFX30qSwg2BSYgnZk2bGV
AP6jNcxtuiUbnYXStqpqCZajBVP+PPc2Qbd0JetBuuhve45G/Aa1hwVkeQ70MX525CbzzPa22G9s
KYeuYunrr5JIUfzIz5Q5dR57eb5jvM5O/Y7HjOGxrkfbq+noBu9f0n5OFMCIrWsAXe77xFgIf0Jf
E2eT2wt7M1ffcUbvfzyFZr9w+wT4H3tP1Ls93Sn2hPm2xshdKdzgeGoFBic+mvfsiKXnJ4wz19oV
v0r3sKzVdYc/VGYLi3pkyVagJ+uAZIywMpFapGjqCunqQ/SYB5pBnV+MsLcWBJXNsnodyj7ScxHp
20ftysDjELhg5mxFuZzlrP7MSJRxI/DeF0+q3kjyhqD4AZz7Y3ZwHRrkbaZJrSeiM+ir2gosCHYA
Q1QKNT0Z8ZymY1E6xT/zBppn6OHvD/uTiI7CUiGMqZ0M+/pV9RD08leYo4ttUCvSDUQRK9lIcumL
7LrS3SnFfCdoCe0OyIEJtEOFDgxrZ7AdnL8YJ8/eLsuW19VGt4Rw1RZOTeUqr/nyaqwYJNkO4jaa
w6odhLFjDO2RZdd6dWWV1OUPjf+8LShYXmiU9Gdoyv7MZiyScGE6msVfYXlehzP/68FHnU6orUWk
XveLJdzbfVHRi+iUL0/q0zCxVsb/pTndEczbLZHptRVHHztMj4RndFvPVSYdC1OwV1aV/5+PCj5K
WC5T/RZTfM0IR/5wIvpNDavnAJpA98lIG7QuBuLSsRa/qYY/lX/ieEWc0u/vAHGS+h3EJ71GZKaq
l14ITuPhoy/S6nyPDikzg8Qoo+cjXmpPfa/ywkZst6qIDmb9Akcj0lYW9GhnDvQVwRxBmK4pLHCO
G9a+aG4VuLzSjmT/3PdXviFcCHx0EzgkH1DjsHqPjgN0InTRnxIfawr+LNGgm5Pv51mPhO+C9zOy
4KPCcNny7FlWkwVE+70p0TAE06cjg939iX67CIMKcsiDH3klZ4zCscZ7IzX7dCm+Ge0pUNGWghiz
Nzg61/VtopasPqlcr3a71jnUZ9zjM/rrRirleDuyAo50rRh+I72CyaBB4LhfyuwfFvyo+W4PcsDs
UrwAgyyiYMOIUMp93o5MdgPTYDXYqf0b6MfOYzbVp3MeOc0YE8Z6s+HYv1RrSTb1etTlqckZagdV
A9pl9dsDKsWaw73+/o3FJulq7JHLW0nzOdC2ddhFOzZQUodV0xmvOCf7YpvCu0rrN0A5d/g1d2nM
c2NXRItQHTBIGvmWn/S0eMv1Jfg6JwlBY/e0dUtbqVTqqJMwX9LgB0moi4RU9jSsh2RYEbMhd1OI
/LKRUOas2fijrtluzni6lzYsW1soXTCptVtt9XVlZCcWE3bc/36u3wCNN26YiXmEYEMQD6ff6MIr
VJopAOW6ezcnWDr5k/EJzOslmR2XVi1D6uHmSpYCry9fjWst6T93rb9bpSW63if+WG8l0rx8pLnt
IkDtIMRD7/AmPJRmZTrAqCGAanNM9qsiGbxpwr+GwYy90kvHJR1OfUvR6QEC7Mc2nwNUv45VfNPn
8YcIUJ/m4fNAiKUgWZSFY3Kmth1o8WlmSjqavxqyHcBe8RafUJeGxi9y0d2o2y9MBZyJIyi7UM+v
8pLin8FTB7lOtnw8X85LH1o5+tEMA3nW7ClfZoHe5L8ovRN5kKAwhCAnYYXvoEEmvUQs0OnNkJXw
tzOf4ds1R4uUri5v/VpDdOzQN7cKMxK5pMMH92u7YYzTNbWSUWWmx96hhPQ7J1QGYPkaAWBCsKJ9
Xq6HpUMS+XGVh5TNWZKQPaXidDxjiGtKdfgLISpfUK6fKf2/uO4xd8MybrBg2e0mwEVZZcUDssdz
fbEN9mDKQW1f0J+Ziohgn/NcwlFhwnP38OF5CnMMZ6+Eomrla9qtYTMfP3yDaeiy0SinjIfvbSbK
i0zzYJfLTHic5w7Q1usACpdaUiqh4DohOC7EKwdWaGPmNguuvgtV9p1lfi+V7aJfgpkQwglQ5nvG
9rvbyTawpDcgozhzQyff9DVa5W/Ka0XFAyYG0VQ2eoRxRMvq8oYdxRqF53hUPk+EpyakVgYLRkzh
8OyjFO356Fc0T2B4ozTrfYVa1hGxfDiWiy9++CJkps2wrqXt739/A85PrISXQdf39Jej7kscRH/q
hfpZliZ5PrwBMzxbcvWu8iYJhYN8QpCZOTfGB0WcwKo7NKDxaML0fCt7dlMn3K3R9DLSDf3yNcmu
aX7FJBw4pKWFbFsKWJLsi3C5eWVGWfXWiZUmC8OD3q2m7/DH1FrwJWwB85j4gsMecoJMoOzs4WFJ
myK0dDCOSv+x02Y+5xyucLasoZey6dnG/c5+aHySEIlVSdGDv1Ky9irh/8/LkxTq+p+UMR1TbHtZ
MOEYC1VcoOT6EyIdRwWk+jOKRX2UbdN+WOrkoHGq1/wxrhns6gPg5Zd2LaIhSIm8AMPUK5aivepd
wNPs68lyzVUyq5vozvOW69s0ChtXwajIoPH9fXAKciEwGKm3FpzCfARNzPaFLGs8FmhNrPzYjNP0
bMNcHWCK7Wlmk3LFU3SGQuax7/oZmjXzPV8T2xTjvbnTUYQ0IjQv0iadCbGEwqbeqn9FdFxQoUhX
2/X5QkJLO2EqEdJCCRmfcn2p1HE8HU6s+LqW6u+jErCCSmZWid4ry+tvhaejQIu5BcxQgQo8MIY0
nGzzb46TFrMhvwWSfF0r1uVSNV2Kq8YB0+QLzeaW1sQrw7ruM7DAYbpKKoJr1h3iJzDfE/hEG6nU
mnuj0F9poiVLZUayGivJ3bdVTXf+ZLIXGITKzS7xUrGQ0/KG+lXC0K+B/cyAQS4ZrXjxQWPHph6H
fjtqSkS/RwgbDa1tWkEYXguXiPk1To3t3Ypza9p+AaODpH+v3Q/hT17K1TtisuApfRm0c6VB5dI1
94XRKUU6TCCqm0wy0Kia4EjFOh9lQG7dDwAnfmi4lSiGGjrr4DRt/vTEm7WlmqDvadmS6cmQPBS9
HRrforxFyZ6aR4QXiZ4r5J9OPxYzALByM63uTGH0Qu0hq154aw8l+kteDUcVmg2+2vqcgBa9vSmu
7AHo2F426+vBxroh4RF+4RJMFw882PxRRYk5QqmunmfMJrFnOaspw8SWRkm7M6XRyyFnFO+W80lv
CcZQMrc3fWP1MKtwfapGG9AfGeT1KblhX9PUWEnZOT8Ilfgjiq8Kwig1ERa9BVPXG6xsYSpSxueh
jYQAH4p1DX9GnAGtaJ/3Spv+AWKCJ5GejM+/Tv0mksquQFy7zsnKQptRdn7QUXzKk62KibtkRXgK
aUztCEQ6KcnTbhnNZsSAZ8LPhhV+sT6TIWj2LuyfYJJGuOI1XfqxWM4YoySq99YjQoJc+fMX1T8N
Vszf+SEeqIA3wzk9oxJAGUE18Goj2H8qOWXtl3+lB8wtYT3OLp85X4HybJtnp0b6m075glmzA06F
AvGL0Us8r+eJxkwZA49lm+ZLAU2NoSknJJjNRfW9ay+/UleEpeg7nSH6ATogQjAMY2RMscGLaFTX
Vk3pu6ytf510u1AUe97IF7/BEX2cB+O4tAtnnyo06V7I16pxdrwV/Ijh7LINk0MF4Qzl56DnBdV1
URe2k+HI96kXfGN0sU5ZsEHVmDieNn7yRseVYcgVKCKBT/HUE7/ZY5mQifHgI93FPR0uipq1kDut
R20DBH2PxMDVEBCcogNApSu2TFC803mU39o5stkQdurUlJno2fhh/7CSE63CTDWthqyafadnxR89
1t/uM5xUGxVjffXpAMyZvK4Ry7Y05JQ34pSxbshFfS3qRMdto0/OErSlVR4hGyBWvHeVb+9kAEQr
ca5Xte8Qt63QVGmahIKaDZlX5pwTk2yzAXHodMtiqCqJQdc2bCvASCGlmARDXZKvK8d2gP3d26aB
F2DKzk+ruxFn4AP6xvP0nElHRhpiY04S9Y04TcIhe4d1LkTsADxX11thCNc55JASmXTdkdeQ1v5t
Hq27f8taLr+4BVFcsOFTiEWA2FO0Qq46Q94xKyl8WczV6wqX36/2lP+tp8Q6lsiHOsT95SQaTsqv
YWZb4Kes4XR7m/4/1lnY3LGPugH8TCUZDPX5Eq6jxr/bVhOVF4o+VKvuGNgm4bsgsjQpSF3Zke5S
3HBslRqGB6Efm63XxdCJQW9z7h7Y+kfALJ91VmLDY3lo7bCTnWkHJL9fEeHdburRLCK9jGqkdVKr
Q5gfsg9uwFulM3TvZBxe1g+sFiLIDjvK7iuis+CZ5VIFVvTyrzVs3v/oq2LrqxXbOKB8GabrB9Bt
tXvdl7QmGZmTfKiOe5UlFhLiqLu41FFhhQnVNyn6dycFm0RQKl3Ycu2BcIrXVxNRTCC0nDXjgwn/
8leAo1KIo+nkgSa5pFzf2xcrc1noSZ1HyfkW451HdgURiUywHQyZs4880jok+MGTPQi2ddI4oqj/
5l2nG+qG/1QQ0SO1qkhoMP0dngkue7bCqiLPNPv1whZEf62d/jP296TOY5bW/givKyCQ6F67NPVq
Rmj9Y0OicyCwRLvNpoemaBLN4lbGAQO+EcQG2Kx4hg8a9R/phEZJ5sIf/440YHw5OJBQkfSY/FQB
4YfRHHwdN1YgfSLHm4xKq85a0Y8cDatOm6pzCj5St+RWiIYySZeFuPhlasmwwr2ABuUSVQ6EPuR7
Y4qLhG+i5Xkh6MxJFbTCG5JXFBXdskXIavS3sZEcAoHOrGkb7kwu7XNbKM12LbB4Bj4zIcZdN7tZ
gilHE3ipW/+PI6n87h4PRt+1rApGk0/8bSXMMJBDLnGpovS39voKfNJCwCcQRpmSp+f1tjk8sttd
XugVJJRPV93d+hAPGEt9nM5q3sgvQZM4aajnX5N9nT08L9viDp6CXjjGF5YIB0J8iEFUgJCEc6aW
5vf5/di42z0mHqq8dbHCdMw4boYfyNhiGsyxYz4bKD8wGdrWCGdSli/J8KyZrV41G6NzF0tjXCyZ
wSKRCUbuo3RKDnAdjJVysQPC6xPN38coisD8vsmiQc9XXS1C5bN97T8fw+LDfz+lKrFTmd5Hk1tO
jUO77JlStdumlgdZ6Kku6B0fsb8c32k81cm7xcb8E1vadqYTxABk5Sc+z8QyMonVtKzCgTm5fV4A
wFeslw9cokMVqT7YPK2Vi43/dpEVPh0bMXEN0gt2Ke3sMr3cWIJw38FMyrm9jsh88gwh+2jap6sF
Hvly6N3fs+ANe1dcHcOz28KmUGyK5yO0C9MZcJ6cY3ksUTaWcZ+acFXsm73mwCqEw2IunAROi3ns
LZIp2/w772bN0z36Th/f8koacxt+GvRKHZqp9cGVIagSz6rUmo9jwweSyLAQqKwj4Z0anGWO4X2P
vD9F8sTg8+kTMsIZayxCdS4BpRUTPmQAh99fjPBylgDUp9UDqG4G4cwvqwX3iACb01nW2Jz9+rHk
3CmDdoqclOvI0veGm043dQI5/yJfeGZdrsHRFNe77B16KBBodF5I6QlKPHrOPf/2awHw1wPqAL4Z
APbw4e4Oid75rGiJPKBnGDEHZKAvHtSxV4jsDhW2/FUeZ6roM43n/ZHPDBI94bFXIXsu8YuOIZJc
vdVpTuh7pdzGS3GkzKCQRiALs7OT8RhYBoLbKgbcOrRYTLSULYWMHWPirOHUFudYYVGstYPOxK2R
qOwJdq4KBhmSrPLQ8F0l+DaPpwXGJ4TISi0som202rFeITLiJdm/5i9C5sM/MRnaNr5E3xLE+W1y
PIwEK5Yr/tTdrgD1jGw1sNRvZ7+3AyCB9xekHHIHJKFPe9HgGOkJyMqj5AvRAcHR/droLxwTUwmT
k8OrDHjbNLhPnzPUfbAuPgELLQ2zj2Hw3oi+B8BWNDu3QQBE0jmkVTs3GapJK27MHlgsKorGB7XW
Zo5pRFp5hhe8dcqX3/VDvFS+rAStY1qGc0BIGwZzxBOrs0FGeQ6Dl+g59IqgfUQnG4f7ElKSR4Bj
GNyFc7OGmolJUQ6JLxb9v6PmOhhJ+Jnke1sXierqAK0m5TvOPodg1w2rRXDoGRO6X0rcS3mTjfYV
ujrLaRWsl1zVcPgvd4TsfVwxGufB9JFeCbVTHSSNlp9jjYVLxaFQvGGMjIM4IHF3LCBNegGjDC1n
N8UzJ2BWFt4WMV1Tu6ahIEcPem7TyjEEcpITH5HXzfeM78JTLBX37uyeKDtNiil35WQnc0rPGdMB
xfpLJMVagKxsX5hVig1gk0y1zr5IVjTBANEkKomNFEcgMZ5khxZXtjHpheKnRjSXK1MNF7sd2FyA
orYSjzO0haViGV+5Xk9+BDCz+UYTYuNTdkcuTsHTbb8opdVXdOj5Co87ricaRjlaNEGJcUfoym9R
p8P988GI+fGBoQh9jkOy//1UwlWFPFwrw1Hnbo5/qvB4AOZ79Xx1EG+0uip4V89Rno8c7cbARY2X
J8kWo3nxwk38cGo4eiTH1Mp7SpGaer8cKPZ/eBFlkDdlzUX4bj7QudgfI4biSe8dQQ7XMsjNcW8E
d5rPej7f+xrdPvW49sYoOWzbAwU7KJbA9GzeBqIw6RqA/FQJKj7UG4EtOIrzVDHFQfsaQ6dgmxEb
X/OEQEzZoyE1yf/pISFZucH2tHsBA4gvudSPOG47vpYIBvu8y+sVxuXcDg2pYSP4yS2ax0prJ/or
0xYGGp8EoxeupISUsEFB5QYHOnMurgfaeEcYkJAZY1jOJdz/splet5IHI/GDe6K/UaurDB1WqCw3
HLwaY3gswjTJ2xc+qvPZmaJT92NJOs1wBxEWvH5SCtdqlljDLVDGop8m8apqP9Gw+Or+cKBAAGp2
6FnQTHebX3kClN7E/FsyqTlSOdJWdH15UswxgGCps42jBF283u0Ed26qnI92kdD9koTjCYidxeTM
lYxB3L1U67ZSfQ08U3iYwq6RqmUDL8s6DrhY+w6fsDBRT+R0aGKH02I46hBkBrBp1y3Lfrzb9ru/
dESI62Sq/o0uYq8ulZI0POmA0h7aeRb1KBu3Chk/BexsmbJ/IwVc1eGETa2NGpEnL1KSHgb9lGhU
Piv/fAKIz1qA8efN/9rue1g7wQeTsiueAG6SVG8Q2MP1bBSnuh/TVKaEkyVCygkk7pr5BJBSh2rD
CEEYsVr91Xcjp2ABSyBa2P+4TJufCnf6AuVFIf7vkj2xsGocHKLrnPIhzXoxPsjzb9Dwl+r5zjlL
Mk9W4W0uKAMAm7MwlokF2avWp5NgGWwsQNRn55/1SDbvID6pTjw3SD2H/pehlIg5kDqa2xswtIsY
Up9DnT4sHvaj8UGg04TJjZ9WKHhrOZXo2T5bqV0mhtspxieuQX9RzkmUpd1fo9ZodmipAkI+M7TN
36pynjVJcn2Q1PyPE81l9GnitsG7F8KnZ8q1a8V1kH4DZKDAcxFyu61LyWWpFoTp9D1r/n4GPWQV
dVqDuyckEHUMUj2FJtwSiJz1H9lwJAcdyM6amKPoBFSS9mMRDLX1diw8IBoj4BVfm40yj3ZoEWpG
0G7O574heAczJ3AAERyTx9K61xmlQrdxmyjFgJwT0n9nM4RYUdmbzymn0RfYrT4vPLEGJB3xrLkm
mxOa0nbU9u55zsLzbxCI1FBrsnsPCqh59WXv4a9bnMCRztLVc2bkY+z52AhwM0SZcxKTtYnUBHuV
XuMxYVw3h9v3yIXUn9WTUVXdACP99w/8JVSDlbsaafc9QNO3LxR1jw6TYHDVFt1wbhyys7OoT0T8
XObt9I9Syo1PA371dXThELivpc0SBtDcVbwtBGjC78foUwQ/cpZ/BiMIxspBrA9cJN9xK05v+D8h
W1Epc1FQcOEoZpgeknGooYO6vpT/ff1eaB0FjIT8smcpb3LgZwRKj9pu+WQylsFqr7vv75ZTmqUd
f1P9YJujwqPKh/qOQHh7pEqmhltFMquap3O0SjjZVKvkEfXuq4niWxSLdYRh6CR2gPqpVIqCzCMH
XvT9XuWnFNySlVc3JYRN8DRGKFATizPJaCxMAA69P5vipZ3YxzrCcTTICz4aIDb4pYF4+ZC1kDGd
LksgGiSZtym3bo9iUx5KDieVai/cR/3gKIf7ST4LjgGgv1VOVzh1niJ0WGI8glb+2ulAE8RPICar
AcPJOSRjKzRd6HJNsz9cvI9LCD6V8n51TPeJxtzZ+Elj2XkV4OjXTEYt8wkSMQ/OiraXB1hGIARR
CTSSJLMAjWhK1CdEOBxKel1PHEC5DglY0T9Po78yhZCvT9BMGuKJ+/Vv8izg8lbsQ3cnXeo9ZCaQ
N4pgi2H5GA74e0Ve3n50Ah9sXbTUjoG21R3Fuyey8Eyizd/XV1yLPakndGFg44m/CCj2h0Dq642A
fR396jKPcI+GR8TNbKW19Y3UR5a3ESnZ26g210E7mVOVJwsqB6sogCdWoXkWJkoXIAIRhewrAQa5
PIpcAtYEepiyEe9d7w44/Vf5glqRW/3IppnbM1HC68Ds4nH75a1RD3bpHI+Ni00bu6AfDrPOewXq
qGtWPm7m58/3fw3lrncrJVwzfvxEohSbPTdxhcAVG3lgMgdlCrBLOwJqT0M/QwX+vHImo5fC68gf
aw9z1Q3uTUG7rG/gf3tr37zR665Jry13LvaaDYH8QiUfHl/Rz6J2K2fuxktDjnLWUNp5pTwdupM+
eWGtTDG29ChFd3R3f5kw61CD/BuRiTRAy23awii2FAALeJRlczdY9sZaIFOKAlFDNHiLVLMMmI+c
5UcXlnKU2LcQ9E62WTf2/jaluwNlG8vsB8RFgjK5ZhVcXoMGYscFv06JFuPXq4GTgdDEN2DdI4S4
xbuR9NXB6xefp6hhkcJ0DPrw4dIPSip9O0rwkrLWVsjazwHPXFz4Y2x1079/3+a1mDBG9yeNzs13
IAfpVw98BqU83RQxXqbZFoyuy9LyAdpZoAF/ZO+mBtGzhwbnSycsJ/BO92S1LkjLsVNEaa//DCSq
VI98Zeo9OYxrH0n25Kazbdo15iKvXvgU15UN1a7B7+uVfHl5TFNQKiZItbGTnYylPRmKN/9xnfby
T0p20kZoamTelta7RO5TLexB6ZRxEybZx/ipHifg0UWclS5fPEut0To62Q1S81qUNxs1yB8AeNAk
bGWLbrbcwFVyu3PzWC/snIrQ9FDnQNKqBj54sQGcoD8+AFlmFtv1ElX3pJwL0iH6kgdtu6KuObAx
VkPR4EIcLeRPuH8g+A0M6lCVHYkPZmqbWuW3QL1Y6kI/JwP+Yd9DthhQ1dY1PP12eYyJTy1sVy4q
CmPBjVPnIcSaHnoJ9VfKYr+EK97URSTs7tQ4kOTzh02tBhAZufen++8/4WW0RauPRFJ9pJG5bSgL
A1LBIKQUcWRVPsnS7Ywjcb1JssVAzVZBwMd47SDXne/ciHsupRtLCmAOhsrWrw8vYkaQzZMM6usi
D4HTuOT+7V5viiBqKevRWi22fXLBSZ6fzMGwhSZnrMm4JhPZLdaOJUtirtJz1N4YNpjldysYu3uL
bdgoA7GAw6omaRhSOjzaKIJh/0ceCk+yrqOyqCFBZT1t1Ve8v84t3ZkajwYSZwvyexK5iXJ1KdwH
IGkblT/eAysqhArX65wjUXF2B5ffySMweqkSQ6xE4y4s9QgdaY+Ob/20ZXXjntx009pJzQuSC7p3
6aBFXGD2okDDp0KAYMLNkUuFgo7fqYbqVW/wOgu0dWJQR9a++FnCUFpTGKRB5PrCm866UlCNroof
DJML9TU7ptNipHVRDMcXIUuggcrEnyJ0hdqc3h/yY4UHeIhZaN35tlF19JVgkKGQzSAfg+vclLsh
dfKS14saWsrFCj2uA+0BiSoxQcG1E1aFupA+xlKmS9qpoAi8CTYsGcqVa3Hq4X/58wQMOIIS+riI
Z6Moo2Cb3vHdiARg8Rw394TsFwPlFxbpggr4Oh5ia+IBIBjVR99Pc34oeDt5Z8J4W149y3P8EL9r
ROhy6yNw/JKog5IxXi+B4FoTTbHr07yUwUL+EJw2Du8bsREwM3UFyYL1K0vi9trZVeym/Ra5CzvK
F/ihDDCl2oUPlHy+UJGJAGzyf3gkz2dSF8TV2H3Nl6mycsrYRDQ1Hx63yvHRsMBz7sIkpoYja99h
x9cSbxzAkiSAKYhMXcwhlg6QM1LviRO49Ey0IL5ZzbMYSgKo2e7TkKRJoPktgJwAicnCIxAn9oAK
OkqlMCWGnBPE2AQBKGYHlSvS+9qT/H3g04Jvxp+oI3q8Oz2ZngRvgELtB3RNyhk0TS/vCddQQLIg
w2AV8B16b2Kze+Qs/ygLXUs+fuITW6reJrFh9O0/dRkSrsTpf0Y4H0AQzDUarb+HESbOUAmB2hol
vH5WhewTZmb2ONkDf+GEKX3VQ9BrFPhd+PlRt6zo0NyxWHFecQqI35ShX+g3uLDqtaA7MXFjFa4s
YNMpYipMcl2R0EuaAkA2TAUB9lifAT1nkuSf/vPIWDnEullNDlmKvO8Zk0LsrSemeKbowz/hFzEy
HwER8ysF6C8Tj54NCdK0ZBDHo4pQvRx7FHOLYSuifbK6ZRYxJYxgLm0pcjCSgYt9SzYTu59nZpuQ
JDVMsnEcJV+tINBv8ae8k3VqzXy20bZ1eIhycKVLzrByWUehIWBs2UurGycX1DR9KyPJcOv29z3y
ZPxjxal7TUiAgXdrCH/32X4CalizjqRXd61yklN5kdOmTNGQS1X73doZnunDvuTESuq5MRP1G+HX
qc7Kt2jqi0uBxZetDT2EOpUSYN+yYSlYwbp52kepQ/ndGdEv8Ab8s+K01wZGOUoJYmbQguPht02t
WMg1V39m5ivuXry97adFpi3FeFEy+WB8AEF2ib7tFOqL/oEp3pweWsZaPUTH4DHWDbidQkLsTK9R
qudSpBdNmdoRFvN6E45s/JqexN0stLOF5ojP2ITp6zNkiRhOCVPqOsCHeQcqia2oxEHzqlwHBTh8
87UWDnTH9LOCxUIIybuSuqwnoMtq0UgTAewEU5B3Op636g0o78WkXPUCDN256zvYwkdA6H/dnU3D
lcDN0HmMiSI+lRsBslHpoSLCM4OOVwlWwzl5VhZJzojKNK63X1Djd4U7Kunygli6k2+XTgM8xGfT
JwRXoxyz1zmKryzIQiEhU0oC66JnKmi77Nt+o74JGK+8XozlqQZrVJEpfDY0Jrq1RpO5p5MAP6Wf
edclq7+pKacnGa4bnYSgawXyAS9pXhZ4oaZU7FDbr0h/IUm/CXlxj28AS6B+DyY2rKEO8KyAyauI
1fut20joDDUBURFRfw6UQRP2ISt3NxST/v8RB4Oq+mSpvTP2WBMAjnMhWVEQCSN6Ne5r/M75uLU0
HdtLD18Rqe8lGxOCL1XB7uXXtGUTbWquk0Etk+blaT0oQLdt2MyfT6mHhTzq508yg0HiYGO+rTeM
1gi8+tHb1HBF0ObYzPDGk5yqIoiC3omrMA2Uvb7Efr/GIYHS1L0RpZZD19QDwIKpr4ZScJ3yyNzI
L2pOK9sM5liTZL01sUbOGKU/+Hx3w5uEJvZ0Y30gWpNnzPVeHejl52P8cSeXdsIRmzsu0vDvfXxD
1OOxnZ1nyQVMaB7/2f7nArR6CRpIDqsKicSLyOjzkKP04TbcndSQzCAsTAgr6R55bCcJsji3qtdB
3licVPItFL7osjRn5ImGn5QXexhx+lu28Wntw+CPJSPykWSkTgjHKJGC5uyq3REbX3lw1tDZg4LE
kllqEV1uTqTigXFezbv+k0JaokquSoMnx8LAGG+5vraR4BgkFALoRe2a2ERPA0ekpL9VHnYSlpaG
uVcBKtb81XUsMUqIoVwc8Xh1JyC0VVKlduLGGeACP+o3HAIr6DiJSY7kydpiSM9cRKyqzYU2Bu+R
q/GmuGDIOI15fqjkMEtKZSgmR8cYLR+LtQcYf0cDmiNSTLTMZkvacXEfazgTUU9Z4wvNDYSu0ubj
tXE3f4AehQ1xevTUgTAy8ybAM8r/uUUEbuWutIlDFh5yRRruy4gCCmymARz+7RIpeeELMRjanp4q
BMry+rWbU5PB60ng38vZjhhKfoSJWJ7aQ5c5xgJvEfVT1fo137R9BP8Ll0HbpfvD8RXA55H0uyX7
B2x/wTaZYMpEEcMOyAYEPOaEGMPRHfPBRtIPVJ0YJGcFTWazpovLsieU8O4iTdcfpmp6RDuUYcow
QQRB4uCcPzjABGdXd+e3JVwIvmoxRnpgp8vAHdTu6oYdwuSsq5xGPPNIJl4imreY3VKFpTy5Uu3o
Iwn6Yc2bLdBxoUb4XU7Lb+hUhx9qYUVGyHqL5SuRGAJdvbnhEM2YBj7Vz4sWOlBNdiPmIf3xHXvi
v30eAnkkj2mQe/zWsCWedFFjQboX+bEtezHsz+UldQb+bfalcnrc4qfKHvXvMXOD2whnswqyLAfy
qPY19GmdF4udf6IpvS7j0okb2f8Txjk/TMr+sdiYU/JDmcdarLzIKN8yIfNg/hv2JGNodnnHeHPK
Ona/kU6pWRqzX0m/EOpWJEWLha2f1qNlF257V+IYfX4LSs6K6LA5SLVuOqWx+IxBKZ93aqDWX3G9
MBpJErDPxJwjl9cOgSCtuUOvJtjWdN92kf0gQMqTD9dfB0CecDNEynx7Eh4iAD643MiDYWpnzFU0
OjRIcdl3WxOKq6I5efGNkTOSfmWpQEeLnffnelrVX/u8iIIWsNd60bXPEbrC0NumMOrjG/m5dKvx
gxE1xZe19VLYNrt2vAv7UnClUqyJgRfk8em2HqvmKT04IcxasfktxpHTrrhiXy6SsH1vmMkue6Jd
7rFr3Ck9v99IlJgUTIUyI3mW8YLY4m03cakyPzgW92AoNMaamFQZankbwLdo7CLCNqclvzg7ofHC
Xnrj8plYd98SxmX5njBx4gRyrfA+VMsQ8OYnp3oYdX4BBG2OrMx8JeT+bhvnsT3T2qJFhOpn5c/v
Ot0BrsuxXsIcHWkO2UZuA4tWdnjvvLZLvSjRoXWuP0nzfQaPihkuC+gPPt6L6FZiRhzySSfnqGGq
m3J10HRNsFL16alXJG48MQJHRbWempErbLlmemfRbON/5dt3gjwBBjGw7QBNFlo6B7MFhnpMs2L4
0HmkZA4SxJD7m7J0lxWpzsbMZMW2eNtsLx58AaoL6KNr4VHrK+2CaQIVHZvim74fNwWa6FtDCVQP
fV0bOfeR08D4odBB4Vwy5nR0SC8Yj90UBDV/cbnIW7ObIW6F4Yvz7e7DUFRGdmVvdIwC6/cTSFlF
M3zHWT0gYzOqXyEp1KOAxUYSFmOlwIjDVmEXPXIm7k2cCuAj7YK5jHc3ZLjKEawmoYxi+5FZAus+
k3U7bwBOId/MQ7l+XMKcbzF10uQEpMIjzMzas88N30FJz3XhAC/UHABN2Qwt1me1dZgJX3/XtKzQ
D4sIcpH1WfehNoAY5wlgf+B1twQs506o7hf+Mt8jCW7XZlp8NShiWjyy9CZvOginhUT5eYJHQcr2
7o/le0G+WCFilfX1t/B4vpQCuRmlqDcrTwEoXIJZXvvXcfq+byCmFGP9bUvmi96A39FZbSWulemn
ywIpuCkvlKAbpR3Rj4o+Lg6n3k53L+Ijj4UM1mkCxsW+kmQX5uG65KEaItCrKu6caRLsEzX5nAH5
MQjDpD2ERWI+E1G4F/dPYpg3MT88zm1q5GfU500QF8XGOyhh2i05o0W4vAKSfXE+lfNYs8wXGbnd
dspntyEsovWIqvnw2r6bhVANIzfhOBV3OoSyeF9Ctj5zImwvNO3jrfAbi+6tlFyLTM//YMnx2K2m
6XXxLozh4qOX8+pKq42TEyjg+53BWTTIvRnkOswQnD5csgv0WdUHcj1vLEPOIk/5j7UMGAEhir9X
ioWbhlyWRzPPBMdl6SQj5S81Ibcsm4zCFec/kWthBFSMoEA+hDFiBmFLtmFgQfHi7lAxuLFTnauo
PJNpXCk/lHjbXq5F/umbKMtI5SNz0GzLVUyfMZIhukjbSN62a3zPd0ltm8M/VmtjoEV4stwlxTCu
HMxx/wh9ACtzn1STlWr1mE866F8AIv7g6+EJH4dIDHmu59bVRe8Ck8bLmUNhgYD2YwZFsczFuHxU
5h7/zdXkwhg4JuW3nVPNI+QYOWeA3xd8RdNh0w9+Gs3GyXXfwC4LHv2MhpGHir182IeImlcEJB/O
6mHWOcT5c7O6kJvwP2KHJSuVHOzq97HAfXXe75YY8CSJNucLDGiOwYdQlcA/QIWaeJ1qFVA/6VJ4
7q+a0lIsxTAaPAC1sQI2nJ+iG92/1o7flJzvU7ZI/dKQOF7PHHshhxVTS1aWgeqtz6z0mVBaZLoj
kM3rWzcqnOjRwdL6FhoNhhPSIMINcY+hSk9yZnnVPy9OujfNZGGU3sYr+vh8tKm0leVP14FmkZFm
pFIDaAGKAcuxf0OjcJDaboqoess2kKjaMjmneWrzS4VvENcVuX2izGDgwYCi5xdg4T8ndVNgzB6j
WU1kVu77NLQMCBV7UWpZE6HvtcDEfGWt6iTvFfd9gjp9CbkyY3Qu2q5qA5lgqNLTXTdSVhJB91cV
VyYE5fsX1lAXe/spQGrcMXIdDVLGz/Pyzy38b4GELEucxOA4W7iEw95G8w4EqzWASXimfMlQgPKK
DeY+BtXiuMikXetfNZBpkHrSP6VM/5tiZHG4oMNtbKMkDlY2T22nrX0UgljCpxp+C5yn1RvPUn/B
LJJoxTW6qBGFc1doChabX+d7qbJVuBb3Ewmi0jJawaFKf0CgpeMTRr0vvshUjQArpT36rre8ODVp
UFtuk87TwF0DoiRciXin2uHTv3Kj59hEFb1o5/bWUOjqt+Qh0UMF/pJFk7jHUpVA/ALz5YpmlDDK
kyVjdb0RRRf/cA/nAeEgTSsY2eMteR+5zJckhfyW/gLtg0+tScqMamdrPsxoWc1+FFlNx8M6UOvG
BYOkj8ZFjvyCfbWrzGb8jOyYX6AlkD+1RaGCL8kTDfd2/NsEFujF5+zuRhbsFOhAK31XNpElfdVr
wgYN/OIxbATXDFZz+mab0L0fEZe0cKWTTxDGK7P0iqSorIjczJG90WvwcIdys9RDWNmZ8yTzu3r9
XKB7NZwJoitiq4eeUL4fc3p+4g28qV9MVH4UTMzY4MuJWK2BzNuevJ8Yvmhsm3RWUrtr08KS3SIf
Zq/QLxkQjdQ0l6/Qd+5h2fWXhV1pKu9VE5OgZaAF/YYnoNDVJZwUDlvgKmR575jVbiCsvmR6LxA0
v8w2Cc3TD28RzM+RM8AITFaetninJuPvhJTdmDdC+/QLnchD2+tivYLDPxOFVoFY1dn3sudFjRe6
XkH9t71lF4R0cxqmlsULVhdA2qTy1V7CUB375DIcFr9iOpV8h2pvEVH0f5j0EckSPxILtMN6UwBO
vsSVKFyifh8zqZ9Ko4qQ8CRb7q9MQBbDDtgT1bHsclg1GpP62yJvnNP3G/ULHJmK5sKW6ymJVdj2
cWlsmxc0JACA3j+96W2G6KuJsdfG2J6ltX5Ahi7ggjTINQ3wPkWtj2Yjn0iekoKCFBuzhPyi2h7c
nEMICM9nctRbXT7IrBH+fctzyP8YtJ3YZhtga0E5Tth8eUBQ6A6IQLqLtZRSE5ZHdsRosIz+N/Zf
81x4Qxfc3MVwHGxsTBM9iB7RGNRkXECz4VBQnUXu9CnwFNm1POWPq8bHvL1sadmaR7J/E8vrizFH
FA0Re7poTyEIX7AfPGuT0gYVNcBYYaRzc04LoFu7S3zysDpJ7+Loah7iy12jXNEgZuelrT/4+C55
XXeb8DMP0RgiyAeqrX6pvBC/7Sre1GF2s9aXpvvt3EP2L/NzyNQaTWBSQkOLEpm4Y3cWpWyWugUH
jUU4ue4vAx1jLtCpusA1AZwK1fTsKLDWJvshFL2qEHdHqKd3h3eoOpZRi7hKw2TH/PWbYD4LAveu
r+4bafzlRc0k1RR5yslsggMBWPumEBygnU3ssjD25sFfdFfX2sjhKLkKrmqO+j3pQRXmm4iW/ILC
emiM7p4EfCaHU9CLa8XzR9MtIuarz0sSelxNrNjstS98hfprq9NRD0HIVBtb3GHjCXFwNXo5ZBqv
43Erm7Ep2cHKsKOxPewWuYyGcArTBSnoHraUFTs4BOsz5QQ3DFJz+gTx5pG2kEerg4QRCXHLPuyT
yq1qVzPkfY11OOWCFQR7n5GAT2Qtn2uQtFS4sP1SjpCfsonVcG8NDats/qs4/wZu2xIXiz1qeDaI
9/YVpLkZj9QRj9S2X8wOuVcV/rnBN2Q6MKQHSmvNW8IR3oQ99aBTfoHe4eZGutJOtDrDSTgXebUY
IlAhlxw8KLaczOOBH8nQ4bnuihj4mnqZYoAKTsd/pjIGaPolTuIc3Dup0h7kNbFqizuao91wjhYa
df8qITb6+irZwvsXk1Biee5GnRTL93C4F8EGkWGOIhkl8H10QzsNUMFbBhmm+VrU9gKcLBHacqRv
puVw66H2sp9eskHtolOXaQb9Leqf3/ibSIxuuW+m+8S5DQTG7zx30oMXPXxQIhU043M02hOmWbQm
AMRCKtgvTSSIkscxDhPkBDFw/MV9IazXCHJV9Fp/+1akhOd5HJxu4UQqaClkubxYWMIKaIZXUyCh
L6OGMF/go3E1ni/qjv40CEOYzw1Vj2ROkbN0frm3CH0+mSto18+Et/r5rhg4iw902vvAv3dUzDlo
v6aun5SgmCxjqNqF+78ha/eNW53oKX49ZHvK7JQiH2yIdhe8o9Pvbtl0Q5Txot+dLH3ZiGFf+NZW
HfH666oF/JgLcnSFW6vpQoaQGA3VaN6A0j7KJ5lWE84C7g0taP6/5BjrqnC+7pfudCS6F6MmojqV
aDb3o/yMuBP4xM7reOshh0b8kIwk/g5SJO9t2JLdFP3bG2mcL2BALCBtiGftLKhFkBioYUSbhRdE
qzUaJnAkY+4/+rl3YC9LGdNyO3/UGXsNIJbiINcGwXjwUcp+/NndHby8gl6JjaSnSTXdNsxuvgMG
R1xM1ta6uHmU9rSgz31d/me5siSwPptIHc9VSkvu3aKKEgQ9UF6+joY7gxiIKjsH+SQvROdi5PAy
F5EsQk2x3SP2KigoU9ua5xQpaAGIQwxRUNOX5wR/M/+m3Ds38uLUJSabgFEKgsBHvbnD6eXDcDfn
C9bLebXq1E8mmDLvQRk2YVq8B4a2+EXIIlk4SP05fUXD3oBvk3j8cgMqVFUuij+nZKDuy5NDpxJ5
0iDJT7ZMuzzAmG2neg06PfNg4IF/ivJSfu3iaRBJEGEzctnwgntvNT8NtTEo8Ig5Ul3aUW+4Ie1C
dDnjidt6mP058S8AFeV0zSdR4LN7xLQE9zJKGfDtr+FjuC71dfvvL6Z+GOFrOYyRsFkMrtAwddkF
EwnsO+J0xQXbwAoc25sbesA3h3ot+UGLBlUfgODHyqrr23qetCVcbK9gmi8ji0IgoSLuLmpsgBw8
cw2q5byzjlpUe/8OyPnOFgc8FMnfu6ppeDAuijY5Mu/j0ihBSLIv4dzVvXaBFZYeCSTLdMRi3izs
pCx9ux8ZAhbZJ5Q1drlSKwMYf4tS+/nHLKXD9OFiBip62lEbIC51UixC5u9VYI7DG9GMf3Cxaiyq
TYhvZMioI/74pycNJScW67uRgPs42pYsQUaCxg73urJcvueWSrN7RzwU3Er5fw2nfg/uaXPlQSe3
1+BRBOAhMw57XLIkQ+J2+0rD6JM3aQbk+Fa1LFRMImS+t6sJmvyDT4zV3uKUJryWBGrc/uWEFimK
OjsA6tosCKDWc3gjZU+ohZ/9pfFSsDhQNGiXtrQ3Eo/r1ZLdpdmjYJyqPDuynkeNRk3LkSDBZNnY
JQhEcL5jBmtHqN5hJVEX5oeZQmGJoCBKJGHQ1QbmifoWeKiBjOkRJnrAG7ZXymRzYcVXafbKKkDI
DxC2JDbzsMp4HIUM3NZmBtf4KzBWON3HwkCNzmaEHrwfXEGo398VlFFoE8ES3CWrJ3fX8mrINgjS
Oj1KPWaMZaf4sUSd+dpqtU5TL4ii66AZW+D0LKuNBnihVPohdYHixE4zHU7EJNsAiUFRQ9L+Fqk5
G9XVK5HJCKE5QXAprNPW33r1WC1QZ+qYIxiuhd9hxyIOF6vteizej1oHXb0qaiKAia+XUdTpoy9Z
GCgbnGkBYp2dCYgtv1o8Q/me0Z7VYlG7hgSAcfsdKyVe7nWQnlkgEKvwOwRSE2gc0b74JH01E3ee
yNnSZrvJ0L1s+OAtSItTb7JmtUiPhmMfbzx3WNQn3avbOpusuDneNFBWBSN+5IAg3ebzQqLr550s
uod4e/CKCkB7wPsJn+OzzNovuOssUWSzKHRG7ETmST50a+qWAUtyd8p5ZAAYzPrnQ7LMs4b+gd9p
LjMs2eMSjUISAeLLb7ghvtT6quI8ysWjLnxKLCcfAhNIvrL7q2jaw2OhIjyTTSH87NiF666LdBUN
gerjZbzjEY0ShvHxi7Lw7cFfJOCev77J8+HrfMy9G4izrLwd2O+qxYpjssUx//sNqNH5Zp4YBLr6
tXiHL5qp/dWgn0dzl0FK7lYKeB9Y8piuYKBUiK1U2TJpfUIZxwPHAVVxv9zmqhAHGIckIgTy0dhB
bQxXmNoac6zuf+QjtNmBaphuCX1hLp85TufHIZ9SCVbynN17K9319Zwq6rCWFcDe4ULaz5eCRekC
Xi5fA3svU8l93cdUt8+EPsCK25NObYS22JAU4EaqFMgGsfJi5ThdrAGUCcubpulbWlj5O2sfo/9g
uHH3LUYka2LFMM0iDI4nW6wYd0sLdlRsncVWDWs2LAagk9WEO34DIvt2Yi3QJPQp1kWeg1gPGYkx
82BoWsgJiSmhchbZ/XDwAvBm0PryLe2sPAUZPHqnJCj0WKvt3YBmlZOviYtUIhib6uJhf8mfDkjQ
VV65fz1zztCeMz6p51AFqa6F8og2HHR6Et18iEBAqiSxWUlxNdzatoN0NqVFhO+cXTWSKnraM+mU
G+AWXBdPV6rTz1kiHs2itqbpBGftJILF99HHyai0flnGBkDJxg/ScxsTUCTZdyLtOglA8IpPJ0Sx
sttpySP2rDtAgFkCMmMqONa6aSpcmEppwuzoGLaeJTEKtSy5PV7BISO+4gQ6mc1I6ALmoROB4tdy
BWoqxejYJPzw69dYZRg1uLffw1YFvGvgU2p+7IQ1h63nBRXLMWkeMEKYS2qrW9O+IcWI6opSzWxi
KZsxr4292d4JFW+Lk78x/W+E1pE8hlm2alGmzpUu0HGSv9Ty56/PLf8KpFnIHD6BtJnngsrQH7W3
LVIWJ2zHYoTlrfIKGglPJMA4cLjChEmaShs6iWxoENiHz4rlHKUBJzspT/Jyw/yljUreYW3YaW92
qt0ynRY9qSmmLqKnrcrygTPxwfn+5DCID9mwNMwdH17LQ9ThTq0bk6W76DoszFZoY5T0Ysx1NvhD
20xm17TwqQ0M0cOEErZ2IhiUqOsPw+uoxMC4BhpuHdm7aaxLBvlhzeo4coc+U4ba647qMffqmOl6
YL1tPB0WmFW2BcWbdE0wXUO/taEG41IXi8V4NX0EBbp+QxM2Y/QPvaT7aaZHubnvVej4tWlKFPIk
3PFcUrHfdTYmkBJrOS/8XK5r6fzB5iRGawx7mw7ru9j9bct2vmhnWQq6RcQNeIaGroYk96YeWbkj
SM6ueDEDtlbz1OQZ2sMOygLe1Hirc0Ze/oJUbgBe0e4wUdjUWJnGdGqR5nC3Sh1qJsy8GibciLH+
1TRt5c+BVZ2uqlTanewd717hT2Nx2sqweUYxHRv75aA+KR8sO14iey7LC8YgVxATfTvYh7PONqXI
1Ta3RCb91/6/pYTzQYM0jcvbFJ9eDj9nqCBEsTQ9hFXJ6wpWu5fzCj3kNdUBFxU6tKhLWapXVtMX
9VunNeZmd1l4Ce6bYRS6f2S6OLip67fsGWqIzN5xSvbIXTUW6R2AWzo73VydsBU5Kjmjti7bykA2
WQvIOS5bdoJJikwQuDCcRW41eW+ZJHj6qmMsnS2TawX5xtMyaVMKOUedwgfSiX7vyMfRaRkVg90Q
k+6WTmk+mopqh5M/E0amKtM1aFi++dYURIE/zkuYvGBN3J8rtMIDFW+Oa8N1YIRmYy7c/sPPmcYM
UJIH0O2JFOHadcEe6C3yjr58IvaoyYHwedSB3+Pia1DBnUD3fa/Fm1MBGNg5Hr5UBlqh5saxtNtF
9UU+XuIkNVp3pew2jdrwMEh4+Z+F0aoic7SBBG4qfF/usgUU5bJJrIqUyQbyFGaMKPHk68QWe81c
JOEOO4VLLuSotjZ3J4ZHptmwSsHaDX0j1KBBiQashkmsfge5AVgVDLi6U3DpTndUOLbnsMoqN1+Z
7h/EGdtX7mJKT9ksHbjW5vi4WdFgcd13WI8R2Zs0G16/mg1hSYJtHWyDynqh5CR5+zVlPRFzqzL7
F73wJgagGT6PygzZD7Ayisz7it7dhjbEfLWrLKwvm2DXvU22ZXCJL29FVHWjv2XgV9Pg0TnUE/H8
evv/mJFHQd1NKLuBZ39WL+RMrcnVTm++dq7BRW6mosIMpTi4Ctu3Xqb11BF3w8K4mqFeGRzG1ZX7
IehgAUpO49jjBREOYL3B/yIziiPZYXBhEBLYOjgD4lVxdsU/nCwvThxddBF7uvWW6mnZNSWGOJpf
wyk1ZioLI8+nBD9MpyW99nF+CoBmLj8wfIKwFGFXt/rCR6nl4E2MZZ12OfhAY8bBaFLpnERp60S+
fY/OlbJ3mbK82OkJh7XOOnAcg6OyFhnVI5/hlExbjGWHXArYdS4hWZusndiT3cZurIIbaTorMVXu
QrIgiJaBG3ASX5OMG5c2rwwO1LVL1Wi9cW9qHWRx87BqRDJslxnyQq8jBw8P7rLbXej9Kfbzg0Xc
/I14eDHJARjQD1zxLwVOy6cjvXAdfY6xNCfR69Y4soD2kw+n9OCyZRpaht5WRV8oQmkEWa0kgrPk
00nIev461p733EQCPOWCxv64wvPPYfE8YXp4dLMDsnqNHcENLxG7scEkbWUTzCTpBpwjsNfo6gs7
JZSIacXBHXrpSzL4C1YAL8mP+I2aRk/HIqf6GutgZMiwzz+hzs2+FSXPAB8nGdqMAbecec1hlxEI
NeDK7yUoHnxAkYZ9fhB4QfZwBZAjK4aLczVaO0x3dKON3Zj5Fo8F+j67Y0Rv6CSylvR3TvRr2bge
BcT7/TnSkXp5YyVHyBMHxjymfOaKeV4cRm1jchUxU30Mw5xZxKcCNfHhJOdl/e1z1Fx1RKRr2ZBw
JRvJEpMi/A7O/4T/XZ480PppF9zgMIhVTPA0MhejQ3BmgrlR7VZEuCUqkhbTzr2mGSOGyrwkE4O9
IhE0BjC50CVt1uVuNfU/6u9GblEnBN1kfL2GbvQoiRMhps3Sa1FMXfYwF/BVWr0p41e0blox86ch
CU0AkVWCyeSNyJlKS7r+/VB5jjGnxSBG2kjhYuU/3KAnjEC09BrpnYM/jBE+PTF9SDPPS/1foear
EH22frF/o0dK5qL2S5OxbIlVjn8qHHyDZpacabeB92XIxsdl1elzU0t5hcmlXCQK64BRfI3UgXNo
8DINXSfoYSq2UPz+AZbSe+Ns+y8/cOxlGIrk4l9gGIQjYwZo1AfEX3SGlL4AJlE+Zsvvrmu28+W8
u++G4GuO4MNVBvyYcbqvDk31uajyebPS1aEZwcixBXCckjWd6BAWuEo+nsT1u/E5MXwL+wl+zDGd
Rez/VojFCBx+g+IzuV+7FjrH4RgEzoLNE8hcn5hKr+65CK6mV75Z/3+jukXH6MIPa9+c7N05CZbX
snEUrJRrHZWT5nGjKbdXRerc5QPGT2xTEy4x6o+v2BcrgiUp4BrYq3ZXaL/154pMK73zVzq3dKQD
cplwy0sPFoch9hNbzS4q0EJj8PGtEzBkwFKZOplg30M3SXHYb/uO5eJIIRIO1w0t5q6+D7IjlcPw
kel1u/9jByeHjg9M3knfIVNFZ5h7L+I9q10CFxEnEKxuTRTsiQPa4AWFQbauiT07ADwsDdJgsp3h
59EKO+rmGDrFJBEkwHRMFBM/ZGxA34zXWURcOPHNHIHcN4exkZhZRlvR2y5rAj1k1bEc351wTfwh
3POUYD/WMFVCJpdvDo3TssBsWx4kZ4nB6nn1S/gNFAmmy5c1km8tSK/qjQ9/X2t/qdYw5jb8HgX/
vhXxVbp4WrzHCojsPOF+DaTHrIKzvIALWhVqCBuCFEGp46rZQmQTsW2B+65fI2SjYAQJ6cqzSN5U
c0UBzV8c1bzWv2Pdga0d8XdQe52CN3SKD4hVP6T4amuQtjKq4QEgO6KHfSMMuLlv34UUCRh09uGp
WshtyyfRzNTCPp6Oz0c+Kp+VPJPVtkBCbKrpdpce4FpIaBoVsmO5+aNTF0qAEioKil5yEe/nZ5EC
5l1scakEVwETl81RJhDty/S3KFeQJf5n0hVFEDmMQYm/++SRde0A21YQxPn/7aUf7yLgwz3kJAFb
uDiniJVvePylVSdXfCSHrooqOHQQ8udf6gbGPzJHaABKFzp26bP91S6ppND59eZtHJ2zgiVi1AfE
e9k8NwRWcEF+d/AUBfXOvpaBVqyCw11Rhd5f5Ar1UJfmnrajOioW3WpFXvWkhNn2Z85HV49C6qMn
Kif2ufTdjDi1AwVEUDI2iz360GYf/RkWdBdgzpyg1140aDrmId6kKkABaT/0FG8ptjT77JLAK0A1
Iv3XZpL6EBgaJ5y/wyqKOpdqYpdzLsxDpyQcsyKuBfoqM9rfROUqfZNgdcorkiOiph0Mr5Ctpl0a
Zg2udvOliiJYmLk3Xs0xwvUlcpoRtXhHaKP1esFFxpniBINStf2smaTPNdrCpSOOb97ow+7D+MOI
TnTv2oGIbRcYHNwgz532sR/4WwtZsX0OpKP6HJS7Ig/p7x2moM5RXuIDY+2UJVHcPRyKRqFOEsR3
l/ohSgWlpAuYy195/o9q9oAKTTuttcbcfPxQdSsBJFp30cgkbaSZBEWgbTbQCWHEPuEPrV4StKad
UfXSoSkdMbHsHiruab/1dY7vY/FWCs226S5iORjO2j7WKFF6WoKXtDfe0+/mW2tZ8DllGouBJKPb
VgolyZjpiq/8FtT71UEH459avGBATAiPgMa3IN6pa0TKzjPc34pIQOf67qugvHfNauCYqgl/kjd4
wvFiycdrAiK3BIYsjhqI9CLTw2CqzF3LMRTuIvDJPXcqE6T0KEe5HfMDDbOnt/mLVMWJtFRsBTqX
pqaLYrQTwoEDcZxrBh0lAQEEhmWSsaBUQnnJpPLPyArGY7cZukTQ08zvxptcOE2PPYo8vxeYwlPk
NvzdmlGy6xckMZApqyK7tMRoKRya+jnZcokxAF0hh6I+CkqIvsVZvHgtFVqpZMBhCzPw0w8yHFct
9FFyAMbk5I6rcJtWUboi32BLMbL9jazHK39k6ev67+0ZkvDisrjOFd6oCrsWgJ0hVbvH1PBS+LS+
np0LeR+EbdRLRhZE2fmS+SaaZlcHQrkgB17mKpiPmQIbJxGiNWx2uD1I8ejvp2y8zkFXITp/nPj/
H9fgRLi8b2dwcvV/k3TXs9KSyOt6R3CYGSaGeFbQDMcfhZ2TjpWgD2qd8BloPVg9rpkjI+xzpAL8
CGzyeZLF7n+nxCEl6W91GlBljkfktebDOr2owhA7FagUcmlVqxgFNnl6QDRQnprdYHfXjzJeupql
SsPPLHI+JO2pab0zxRJLoIxAOcaQw7ItxOvro93tdOSqhMoDL2Uo2NwDlw9tjpz4LatAl3HQPUVx
jgCizz3oTpXC9FHFV+wr7GopbFukqHkjXT0hFGyO7pMx7DsBwqvxPphLxaWLgy7wkSvQfBV/gWlf
zkziJNWbVTPisPIZjRnad+2az3F7htsrsDY58UBWjyyPhWssZdHr13Db0OFyfVRn8b84UKwcvyn3
YtI3smljA+CYKanfWTjhi21MIoT8LX8rWTC5MRdfx0JpwMM4d36Tlrec9eR08JkvOFwzZlLLcY4f
wBi02ztmbBs/IDjVyJb+uDgIv53/8Z38RFHoK1NSi7u5V9x8snhttc8U64I1ROip0jfaGJoE6lBr
hz/1dOQH2tvT4pQjeM7B3WO4uup3YybR+L9U/lWUB523zwET5RpH8F+DBSTufow7OadgXYxRkrcu
Ct3gk8RbJrmbvKuLHeacSweoBE0JTXSbr5iqMCrU7s4vx21D/nR3MDDIcNUOO2XPxGLhlYTqs+vx
mwilZCzsGdC+81CZVrt5T8jUIAeLk0OiImrSM8HHmPAnqEJaoSSjgWP3ke21apwSEme5Lp+knUSW
n7EC/cZcdAkHNy/vD/SgHoLEHW8RsIcPXRQROoZQw6pxgC8gwEgragcdL57EfJMEICd4FKsyJWda
TgvMzhQDVwykpE0rjFcqhk30sqQivZfU153MFrpu/w/2o9fwH47AE8rAy72XOApfVQWAvRmAanst
GNnP0kgRD88/R/LcV9wbpZwoWSrG8LKMIWohESddUGq41qI1VLX+IbkU3ktQCd5nLzfFWR6D69Mi
czZOC1QBRSwNWIs6UEKm5M6E0XBvFxCuOp5+y3E9QYLZKCK04WQGzc0f67sWtXyWcpnS5bkv0cvt
HP8w7eGqkO3kiPrTViE9Uwi9X9PveaQ097VhWUj/CsFH9DHCkP+coJixuNIgNOR1G7wL9+kmm2sz
/qEmsbr7c5Jiw7rD10FkRcjyj0VWvJXVlb/PiSy1VIOIr3NicSY0GDy6ei1uCPEK1uWSOTt19dPm
4U7veHJhxGzjnaLTGCDwbdIk2NY3Zo72QMsp5R87KFnj7UdyJ8+4wPMl4M/DbGW33Xs6vDRRt+8s
uaFrXOoskZBafdmVUK05hXio70r38z6p87ubxVzTXBIAAWtBktRKsyPvkABAbSG4G5Aye8pVz4kk
saDJA7v4soa1zgx8Lj6gZJASUC9NGguUshZkLdNcMZ779zsvIpxayNDpW6ppjuh4tiqJyA/njOk1
nSi3EsBVN+V6arfEL3Vn5m6s17hAAkW13fzpWX41IJgYbouhr+ZGrptEVaEmV9hpBoT008SP4bUQ
v3IDSmqDgrnqp8kzUZ5/kYcAhRRLl7ycXs3Pe/IDOsc1CD3OLKvKvXfT/yT/u+SLa1sltTB+o7qv
X0suGKfn4N3KoIzFvGwlj276jgN1ybdTy520NpgS2CprPg4CyyR5CRggVWbFVdy8qLfhB4rXDWdQ
HVFwFS65mbnS8QmWDCCnRVycw2Umf57nLXYW6Wam4bDmN/ycsGlYIRjp+XktOgkdaYRPYB9vjgUN
RcFiBHKxIzUS9X11nBlysmugmTaL/wNW0MK3UAdGvFmmeuHhmUifP7Q9VIQUk58bOO6/S6ixru8p
CFwnujMS5K7pZ3McZ5+LCO0fV40AZL504d6v1KjG4WUwrNjjkWgKREweo9qsuGVXqsIU4WxKo9fX
/wymxxqw6EZDMF981tz5syQULISxRx769wshx+kgFPd5EuDMYKiMtpuuLsv32ZIfTPcGWkthAQsX
MqvTj/AtmNKI570X7g1vT3UTV3UMGFAoPB29b8n0YDRdHiFOWY93Q1+ZgeqHWR5lO9PgwvKHhvzA
skd03w9jIXM0rstXrYEH22AnD4W2yOJagEBX8r/oSjW32OAuqecSs0k8io7l8iwGTTeD7nmvYyHN
c3yJ5ouX8lWK/L7Jbk3SeO6OIjfwAA9uL49XPwHBQ1p17OqY0fQ1NuYt5Fx85Xyw9ZPrjoSbYf7q
LkYZ5VBIhRNDssYox10jodl0LCTSP4xMjv152QIHgwob/HChwILsOl/s2MCOdc3wR9OLMhrQLz3H
mz6zH+ubzz2s1EjJ0AKd/G+bFDxA3rsjidySTUZ75kF5vW9WckQ+NwUCg+LGLPOsOWZ79MLSLhlr
ydQY+fNi/wieaJkgHdqVsEwZoswW9gf/pBU5Sc2jH0H5CawGP3jFMVeF75E66JdP8wtcKpTDcdiV
eepsp+tllBbiSd7TbWhfdDDgxlsxkj9jCktVejZAF4EE9EZAXeD0XAkPT45Vmm5v9isaGms7QI8J
u3MlXNtEkrqkbdrjqEU8ZEbp6l9gRT7eE8O2ntYUdbqM/7EFGjuXahAN1Od5PnSICfl2uts0aguY
K2T1AyU4l6EnbexqISh3Gxxmmf/AP1oVZRm7u3Z07Aiy8wmYEhhJhYStSFrlo5fOozvM2iuyR2oS
DFKzZo+6rvlrdCG8mbQYV/QbrzIlOo+hmmuTd3od8diwsuCog5GwLAp+5BwOQ5iOkkd+QiKZq4x6
YnTI0WzFujEkgltjmgjhmp4Azo4IenrEQURzzqVDUKwq3AKqk8FnwE5k3Akq/iMTrg+AorSgT8i2
7fvOlvzuF/4Q1uOYS8GGdE/jDPiJOCWdETlSM3NQpQ0u53RINEAdiO7cDoIjvpNGas/bbtIEJ/U2
eCn3ni3RYQzTllJndfkLtdzHU5WEl2jIkMs8iiApD/4MmhpkVS+d77ghAlIXJ2c3GRiRzhvhfHWV
tGx2CtwD7W6X5p7smgPoLXMkDbut8sd9SuyzLdsTnCPj6OAygVPrZO9IeL39z1VAr2bzFpRghTac
F1nPOMQ/9O/kRyjfHQbQU7WtZJQdWivoLxAS3qMnUXx0SaDX5LqQ6WjdyJMGNey940/W2kEguP5H
4u3FGM3IPMGn0c0qX1djvsI9UNKoi30PrAiNNa4Uk47WklYTtlAYOscnPK+fUkWZjJJPaUaI9wr/
y6TNZDsQrVE2SGkoCSHah6RdZWUZ1A7U6Bo/ECgPafDWGCNbUR6qCU4lWXdmzqD+ZgagXIdIVarp
GPl4PoDIhqzeH1cDEvzujIoGkUL187I7KnwRwrxWEa2EOxSSu3wbEqZivGVP9dTbL/ZWvDl2BPsJ
CgoT5PgAoWKovI0HuNjLdaXkWMaxkxg13hOOeiekf2vqmBYGW1RdOxAqCA6Ue84SYsDt3mv8utM8
QBuIiplXsehfgW76jQHw8ZjGLZ4e6yUCHvqgExq6MT+yA/3gy+bVl603HRn0nImICIACxBaGu1Rm
Jlav90IsJ+i4EVHcn4R9nW9LDvs8If93DLdyPiPtHq+S0S+aItaY/hQDd8wQc1RZCg9KSkDeZLqg
EmNOYZEFPyzUYvfca+L8C1E8R88aE7hMjT1sqbRt0TzvRswVxZgIaU8H183vq5FgyP86g39sbT54
EmWu+7go+7Vp+k/lwJzuRJgrqNhT8PWxLP/OCVsT1f6epSta2KwbDCtASpFJpuCMEVWBMNwkrvKw
tim9GDUmBAoGcBRmgfoxs9b3NszBk4SZizs6bp10wPS5kd1yCI4bECjBibPYMu1j9kIsj7DK3khn
fZFgcijg1ttguYxf1EbR4/fyunKY09j4b2sLnKM1CblAeD4/9LKIKVgMSrQVJFLEBxJ/DPnpBC48
cLnBKrzKKo9kvOyw16MJwhqT+Q9MQhw3YfWDs81dLVclalm45C6x0ky4PKv3JvZ71UDsk9VLPDEw
5d8dfNLyjuvWLP8SCk+xcgWt1gM0E/5GmNLQvDkhFALCcpAFTOOjxrYf7nNc5a/3LV9HOwDHNa6E
QA5/IVJ1rGHJhNOtQauFlAN6f+A2tKmaJpIDKr85QpfaabNyUUmP5LYuhTRVLtg/4JfjjV7kWEdB
JjF3m749Q+G69cYw8om4gWKM9Sef8xQhiJR3c3YxnQS4or+HgP0R1GWUD44r4WMSFoN697z1PA3w
TGIvqOHhzhLRdt1nsV+VRZ1cslpEV4ffMJ7PyDntj3kOl7gMchz8Ftl6nwYTxJ+T0LVKadmRpxKp
moT29lvuPRQjTIRSyu+DMR6+uRo8XLxBzyd14a9Zl3K2DA//NNB2/Cpwh65Ht5vQvlqRUb7I+ptu
PSqH4lES1URPrmc9SziItDkqOp4sg6OynXnlrI15TJY2+0jIA2LrtS5uS1jViSe3FNAzUbeP4yH2
cDhsw3lNn6AXRHW9owNvQm/5R2YbpYvcEW0nnXr1jv5VGAiN7rfuAH0wckTdkMYwcggtgfQaZVJe
3NOVS/Yc/pKAf2YJdWmji8etcXjwXUji/AJoZi/oB0hMDtgvcvBOXveKERZUYLYqMvpFC/b1EGT+
PauOKaEZIolQHN0b61VYgDrflfee0EDvzrgiUB+E0OpgtU175WT5MTsNAz0KKKhcIK4SjqU20Nk8
Tp5VNPvoJoWHlgyakoSoKFXkMlADJ7p4H/2ge50dliL3eMr50ELZRonEddEYh7ptArBHzNzcESpN
vUYblxiTk6z1qoc/Q+QR9SLUgeYnmbCmhTsU1iilQrT28sTutPr5s5CYK8nNF5bQrLK18uGq9e2P
wlFtOyiClZulL2Q3LgmVud+dtZDJACbZSlVadawyvX6xwagxFdH2o6ss+KB5VmMMXOp61uytvhjr
Otol/0qifLohIwWCGjvqFenL1VVr+cw7p/WV2HMfyGhO1klXRwKb9Ao/Dvs9szHGP/Wl3Mk2DGJw
TXDTkRqIH4CBRncXwxj9rH71BoqRUht2f0iKaJFvNJioX2rrD1MUxn+dupT3M6mqlNA2+s56GNtL
0bbfZOOzT1klnPPt0Xu4dWxbbvcGEs66GRPxTraGMF2A6Z8To7v2g57qCbDYu/V/RK6IBcf7VJjV
IvyCu4GvBrAMFW/1NXt+ymHpcIGLgMO9Kac6ojbVlVDv1wS1HEIGCpL+nLZc2sBRJvrGKhgCHEyB
0vr7RcrJElW/G0bFp2hMoqrOb68rdBALhoJ2o8/q9Jpjp11QBUWUlk8/NWjdHLHUnBG4/Ql7y4Sx
k/pv2DlKgCED7UO/JAA6daYj4Pz5XwhcqlQglXmRtthzDJNpN8c+aYI4T6Mynyuk5ilu4SsG90r3
mCvyETJOrJjrMeYTQKXfkvcGduBIfPsx/szb/wG+PeOFFAZ6PdR/c7NkG9tCz6xKGBJscLKj+C40
axBmSzf0BINwlZmBWgVo/Fmi6RqaCZR0D63HM2SQx166uukfnowMk/RbGp0Ln16rIrFjmpsK3Lhd
7zANClMYzupazxrMdb/+itQt5lLhinpQSJW8NKm/wPOox6BpMoo7jUQ67oVKkUASpmEqRPguhdN5
lbPMtJEegQKFEZeNdqNRfww85r6u3hdybm5IMX9SM4/FySg7zI/JDX/qL1e1L23meaTeCGAHwEZM
I9az9Q5MFG/3zRcDI0H+oiJtl5YJp3j96P73ROX2fZjPzGAoif+qGc5WnEsEvkrexQWNGmr2hDwm
DXCw7aA/TA3lc/Y+bQbTNgSUp5B573k7q+KRekrY38l/g+V2Li6SSOWWI7Dq8ql3S2jJWevyAKqE
FqKeXBsft3YL+SVg+taqnrqXPIb2nECDugsMi619C6PvGcOVF5OIKmCl7ZL3XLPs9tiykbnPuxWS
/f6onQ6XT81/zdONDLuVfn3GyJQd+wfPLqmDtSR6l2UhXG9MXdmcgjqV9QhXfpNkyMIZBk1XSqsH
SHwPVzLtB8l7ZUxix3XsbypxBMd8yRcFYBMBiBr07QtOzGmbO2VY+VIyzZKLsLbw2tghAjNULr6x
4LXpooqUX8VJgZGp7Q3kfwQL8Llv9YvgfptDyAdWsEbC+d0IQoU+uXuUt+gso/O95dQY3v/okfCr
PcHNi7zkV8uJ4PRz0gr3uTZJzD2mEbmd9gA5QsVEV9BHFyLoOdXvKgAzMjd+Ydf6QVA9oRXKBBoT
N8Rq2Xls+TVKxm0nmBOqHFv6RlAl000Zj8ZMwSDYQbmcylEJtAX0bB9S1I/AkoPLgXfD8SuY6vDf
jHYkTDjvIT3+2OJTagDnu/Y15dby6ceTSq4kwSOG95pHRsnKOz9a+dt7NRyFL2T+s9++p50zhjqc
ZxJPy5Io+MsHiKW9nHM4uf4a5dN98vqz+XPzwWRRbMHajCHRgzGO2i3yXT0+f8uKW1MZZ72dwbTE
k1nL0AhjgTVQHaq4QnbPmkV0M5UVOCaIaSDnzjdZhA702+EmBrgTYcUPiC5WLwFn2Ox6a8qajMXl
FBfK2/ZSkF2JGstWdaDqA74xdtSzfbhlspXivKo2KgeNuASDzljW0k7FNp+BcpmfggNNq3V9a81t
x3V4qk5Bcilzq30MXyDKyiHgv9VVCcAP1wPmC8A45+7oa+JrxgL/ENVDXXNv3Iu5Bft1m4q42Msk
AEYAPmAUgEscNqrjusizor+qTGskyKfkEfVv9bE+nxAmsKSW308J7UBqnTXe3dxlp7dDm4Trao2N
jCZK6gYh0rm01lHqXOZCxBBHBchGvwFd8VczfoLarTlY7PZi+RpMXO84kd0gDFgzwG2irRWlbNuf
92d+hRLJuqbh7kF3oaDg+MSPGmuCULD34u7fid2RnD1sDnVBAVxJuAr7s6Yusk531ymK55JTGyaK
TgC1t9TZ687yKq6SyQ+EQMrtpZOvE4vxjVxfeZnMCqmkE486frUQhwtvEvzUHnm6Xu/YKMGn5BdB
UzuJSq8wPwgQB9dU+5aKP+ZuoqlXbw7t8FwyCx5sCfr0oQy1BdCullWSf0sY3yuyX3aZFFjY+Z6d
+P36dmF7o6hHhvYHtmAKlWMwjcp0gmngwGlUIcFvYG6O66bQwkS79CsDTnB8OdfCgM8XbfhdNdZB
NQGiW94j4zv6QqUQvXum4GCi32jOdzoyTitVTkIGxl3PPF/3So6qUUq2E+U8jlNtAb1FnXVjQnKu
mbx9kzHaLuJp4xpUdt+eVq+OVXNPdCBBsNruM7pkx9s/QCrEL05AfE6oo8s5ouTZ9oeoFXpbFWh/
v5v1K5epDY3H65Mmzhl8OBbVGmmkLtDxBvXGSgvinsLCPnF88OHJn9CzYgm5Eu2ZjdUjdkN3Rth+
v57UEYBREuFS7Kul/WZPDQrLCvajQ990mPngpDI0+3KwftbfJgPU+lRy3VHRLqNiib+zsQBeuYoJ
KdORVN3l9KXL0iZ41WMQUESVWT9tO5nLvIaaFQkCTR/j+C1KMJuLv1PnmNSlQzbWPqlktslPvxzF
yUyPMP7iULxNWOS8mpQJOJ7pgtTXYk5Hy1z/Lc8i/FhZLXpFsj63cBak7ukivZEGmQvfeVsPB+Kp
mi5CwmnMdoLluCDuKViGSmAtAzj2JEcRqZKse76FAekx7um32yk6bXvyHAjcUycDJObVhd7S8BzE
udCmTRnumKIYw9QcxroxvZVRjXAQwrojFVgff6aIgAuvJsId29FqKZYb5X36RSYhtwCo5Y/D4ICH
NTgKG7TAnRllGrayYh6BdjrCSUg9j3/xsGEYazUuuYiJuibj4fO9bLhd0g/AZkyGtfhIA65cAPgi
ce6piFKIBZkvF3xNzmMDLJN9JsLq+YROqlg3uBUsNHZgMI6+bCVxuT9enKN+c0Em33yxvSzfP+oh
3OpTH2kKq/v+NLwXGGoYzu6rLt37K1vc2RkIzDQCs0KIE3c/ue+zWi/sKr02FYpxrOOw//BPo1Fo
SWZPYP5evDXZBtUtAeq2Nr1KB8eO/wxLksZAOAiN+QklnyWCzfjv5k5vV3TVWHQjq1eVvcTgbU1c
eQhG6LP74Gf8wT3mGBG1fK28TRDuImSRwFX4s9RLNlo+KFuUFjKMDubz+MfcbZC8nxA8SmkGUeaN
/HqVWSqcttq0fa9fRGpRaK26pKEegdR7jKeohIOkXpASQaKYfND+Aaq7SZ56LAsJJztrbUXFpvaW
MRfOOt5E5no5TxyqRLQaXQuqnysHxfoWIDuhVd0Fobnl1i6avmhkR/qnOxBd1siV5nmA+6Dz2Rb9
HMM2dy+XEeqyt5jEM6Yn30QTwzcO0fqegPgv7zYcTQ8YJXkPdMLXZ/CmYuFioZSr+IcHrVKKivOe
nlqcZLBQaL4rOjFhsEng9MewqnWyvgmTs88ZuHeNZ8nL9X4c3/SrMyQNBvCp7ydnOD4prXr8wobU
9OLubsGht/+PF3f1FV0NS46kWvgfo2ari8yPV73ViZx2G5P5R5gBzKoYJtze0CVafmaLjQtkMWU0
z10qRzLu8sobZ2H94WB+wnLTVx5neth3J7kaZ3/M7LbJIAnDA+XqN0PaE4DGZkKcD/N1PSbvupqY
zgrZowpf81UYJwWhKHBUxm6qWo08S7LdvCSJXte2YZb6E9WoxBDKaQ+A27WfLo9GkCEDkt7b/L29
oqNk+wxnpYgVEy99Ucx5wUu6EX3vYpHpY6GkplsqHr0QJ/Iq8Rcuu5sAhUaLZtCw0C8cqKEzXpUl
mACIVjCq9IhYAEcxCTFLQqVl5xMqM35XTW8+YfRfieh95LEq4jeDLZ4+E9V5cjSMtkdV5Io8w5Ct
jmYAtXHcIgFVTIIXFrvA55XOh2hcVyI6D/OrbeqoxI7S3OY13GC95hTCA94OC6Ovqev7G3Lt+zRp
8KqSWqIIMpjryDeNOAi7JQMYht4GN/Cxoi8ukflmNCQLwGYiDsCnyoYupkyZYCNSTcBvcobDC+wl
nyDXXlenA+SfuwaC6mIQY63SXAAGGzwIT/yF6OfbT5cV/NeKihMftQKO0i/HD0FeEzcagBIjqp81
GCHsSeNudM2XVx/w26/MqMQ0cpXxFYodrBRKC61fMV0PnQMBUanQUKbhb500nFQK5CyLtVydPTYQ
1PNh2mFe3uFgkGW4n0x/tFWejfGBaK4GpyJmRGrv96A/SvjUfBN9Y7bzXdI8zHpOM/5iWzdIP2/V
HXwjGg+jCeseWeL2B3Qnw9e/pxF+ykpKrZFki+jNq/3N8vIWtjXTGx1nlZxxeHKCAar5MU7urG48
enuwuQdkRUqVRAd6YmweHMbkAlreVtATjEa3jIcHo+pk3JU+tGXoSnWgwA6rxxAs4G+8joDLa1bM
o0AxUCfprW/BN1sGsSIMJh5m3lfsYb/cS0zuwPTyh9IRNfXKZH221Hi+OBNunXlD7AdCh47Npv1H
sEZvyL1YftwVMgSzk8qUrT2heT1edIl6UQlawip+pn89+MVQxuqffczHyS98HRaVzGm6O5NBRm+C
l+THovSscRnlkBR0Nl/09UvVgx1FcGKU60pXvwyHhqwFJH+3QVd4LSby3sTlvUCOQTEF2A43li0Y
5PnleNFTMGZ/nQsP/whFjwRFLMxHjsdvXJCKxb5ZZmDYFRIAYs3fZ+GZZ1mvyDwURHQ2jTWkgrSM
tnTD6O9bU3B8h6nYfK27C5lfioXiiwqBvrw2bTjcInkdSN5EK7WdGdvTQCN/0pJM9yWZfNvNMpu8
X+9cog21xwQdvQe8PD6TvUwfV+y9quOLJQ3sdg8pcfzWyNVKuKeGzy4jaNF4rZTpjP5lEF0WAobA
vYiK9Yk7Uvjai5x9LBUGStYnUKiUSYkyZs7N43goqx2oTbmTUWI5FOwxRMCQTiwhKyw8pjbxaJZo
slqlpPnsaMHzKp8a/HPu/IB89P8RrwJUQmtHUGMUvcsonvh8cVzj27JyCF+YfVjuhHvExL0hObJL
rxaXtuGoH5UUJF/Tko6kjyT6xZFq1PWYnXFPt/Lwyjag/Dao2azS476h1LffSbX0vSOPKaeT9gvI
VcFIYMlkYtLdi6CwWtsmX+doHNyNR+piIN/0EYeo21DMnERFULxXIbVVVu6Jb/HcmBd+pewXgSMi
YXFH7nu3c5fTDCpzwz6sw2fH+0JzAernDIN+YGaTiX27FoBI8Z9xAL5+cq5iT9O0zAMXyIzOpxN7
ygV4EvgGfslY+3eVnDhw/6Hr1XHXQjdX5jVprlunqJVY+Z4xHXMUMEHWQVkIW7nk0HrY8IjF/FDz
AiFIxte+OFz2xYU3jp3JX/AJQSErzxA6xbmFTlNEy2Kls07sEExBFdMMNjXwpIEgj62kjdN1ylWo
RdkRtABN2KVrNQdSF03HrCr1JfXkf+vX5T5RXD4eQ2nFEmYx4nlczCyK3R5mEjLysNfPCq3FnBwj
H2ANaPK02E0EtzMsOoawL5l6s8F/C7sjg1npFkKUFZ8jinGBtQIRLVjgn7GOwU3EBVrgqhejp/G5
LRCVjKUjGchEHyR25VnVAOPeduFE/M+oOzmpVTFSoh+0X/FpXtXC0AHeXhOjJEp1eE5A/WQSe4jJ
DUz0rC8kfQTE/9uPGXSw9E4sTbR9zU+whW22YusgBLgFY86NPP6FsSZyMiBJxqcOLNUfqsbIO5s7
HCLPDFmsfGssHInFdmwr0rWH7+YkXiLGJ4P0+WasmDcni9ZufqCjQtfh8ioD7m8+Z89TVzW6lyni
m8pml9ONrXEZSU5YuKOwW+cAmLzQqRnbszG/Vmm8ewYzwFp3Y+cyreipNPqDBlwMsnx48A01tmTj
t93zTwwEpcKaCaopjZk3ai4vriwD3Z9Qvc6nd98fh1goOB/yZTo4KX29aewIok66DOMcPvB9iaUL
y/4MeKjHaz4AqRN8QssajLryORM5y5TW0oPuyc336EKoFmTVQsDQ0pd2o1ELtIgptVdS/L3HKBO5
2omUcTqn3PRtCav++p2UaHC6czEBV+G4yoc4jY2zU23kv1baU7PWZ47dLfOUGAS4peSvRaDYKSPQ
GBMwyw6RtOrkWxnaCpMBjJYxFo791n4efw9BvfnhCjFrU9gQVP7jp5uWVlSEJ+y9kZoFoKCoqfUJ
1ObPK1PKG0hiCTB+aTATLMnzYlPk4ysPnV7CMRoI5TaJwyPJYgLOCUUKmdW6of2uLk4+2Fg/1C49
WuBNEcajbnnDIjjOu+FzkEGfNf9b+T0oqti1zGxNq8b8MNovHxjm7IzX5sDWIGwJYN3YlvXLLMqL
Ib3Zwv2qXIV+nuzT7+U/uXdg5oPqCNMprxyqlSfDru+PdJGvB/h8l7L8G2hZp1yTEQLDeXXWxiiy
71oXJWR0Z7krtl5mRyAQaT53eeOmRjBiT2eXrPyqgokuaGmG5IJXcDQo03+3U0OvCbQKMiFQa3Zz
PjXfwt5oD1JjeGOEn2CUc2QvSs+Ei5SUGeG0ZXZdrtw15IwWZY1Q7IipPQZJdFPT5ue2jvIqJS7J
1C6jydwF4iTMv21tql4qSnQ2hBRy8e8jS4CmA/lAAOgkpFdoBmINKk0oc+7FD3kDG4nJrL7Huamj
1aMLI5ywpCQAFBzdq9C9etsHmyU7WCe0Go9x7Y9zuXPSKJ3GeKJ5PFKkGI8nLhIrF3BnTcg0P+qn
7/5r+vTSGte5SiVqQotG1UI8CttAK4WAvfgzgloz07qtGg1HlAM6AA0GyIH/9epFl+7m4il9NPmG
7a4gpCPH3ZQRhoDU/3Gxy/n27wLN8Pk6NcBtUJc+GzC206cM4YfbJktHUWsvpYEIDHJ1k9O6vgay
jZc9mXo16v7kP/fvLIAAX6421vpe0DnWkmEuCRr3X6rBFMmlf4ujXHBwi2AyWqolRjm4HM8V1N1p
V/pxZc9+fAhgSYPwMFd7VxpTeum3cjjRwNDPr0iYBFFyK+rbnkno1OlUveS9xjs8jFd4DtQNLNyI
FZGixOdBaH2rvgd9bMgbHHWXWb5JRMIXq9Xg3GV23+jKAGwLmuXr8z6CyganfSJkByFZRK/wmTKA
wCIOpOP/GiawHrXOGI/EiWAvuzkACnIwVXsmrOebSPwMID6MiZ4iJGlWiRxQhR8g9NfP+q78biel
NQk/Juc+0C9z+mlYXgpUlZKyjO/MmMjiRtoiMkpZTCORC15zQ5tZ4+MLlWh4461vhEMDOcjy2keX
fIrPkhKh66A42OOThv1PMEXA4mKA9UTAcjXM9zLKugdTVfcvbuKwzgKPbXuM+eV5ZK4cMn2Q5SmJ
sjrodALj2lZpGsNn6ZzeWLmaab1jYEV2FVZsH739SApBu2ftzorhG079Ys6XK2nQTKZVJjQghfEV
ychksFdsayQLpntZmZlHTJsgNfYLTOV1s5ymgaOXUxKxsvPj8k/QwdMPHLc+h0+vxOHgRWt+VZG7
OVVzrqnBfMaoc4GKWG6WsLqXDVHfokR/s8E9+yrzpCLlJanzDtmF8uNJ6jyNB+9KNHzTQY700yRM
jpmhARg8EUCltBnFlhzS0Vx/P3czfD6LhWAUeNwvI5IPlHQsX/BTT5VJHDpg4jGTemDvN0lfY2q6
lI1KHOX+YZla3KYQEN6SHBH3oWRv7i6WSW1YG0ZYdz4/OuG+3FtJTcXEXztDi+xfVrJ5+bFlbnKo
amiGmTtWGkKF6Zq+N1IBGEKpcgJIftjb9tmsxynkRKNyGZDxLRPbc7wmqsduT3T/Sl5VQvxDYyqh
1jxNXpgJVzzGOuepTNBO7HzrxWZZnXrzN/rYCIGKSjOXe0cSApTAILgZO63wJjG1AEGBbO93wMAF
q0jNGGy6xKBPbM8eWiiMnCYqaAcyRJE8MIOgiBgN+oOAlUx8VT5IVEXoIoGX2m6osDgAZ9GDSC3V
p/BufojixCapstnw99vEH4UvPGpRlsPTxf4tvJTkgRwjBjq0X04mkoQILWxVBCAn5DutIpctSPKF
7+vP3tSjoxv7pGs78wVc/e4wPz3A7aa9yN20E4EypQXQ41ZuMLFnlcZr1tvZZrKNtxnZxPRqu1Pe
oqvFNp453Ix2feZEyYPp096arD/3qnsfpdiao9nbxhW/K3sL3pG3Nyc9GqMG5XbXFnXO72SOH/PN
ha9xHq61kUIwH3V3Yj2QEwjn4S8ronc3P4YE6q13otgd2ycdNmD1+kMogRYQYfe+iu1eRGIF6vPx
z9nntWAIXPvUi+gjYzY+dkmerQOCD/SlY0w4wckvlR9/CSWVGPUToHPBjgit/H8G9IhJUvP5ZMdY
5SgUlG83HrpTmSf/prNrIgNa/GJz/PReaSaO1Q1GP1PUtq7kG2TTM2dnrBScRpHVCfN5oUlQcmwt
0B5kEVzi89GJlHYx71isMjlZe4mWIe1rJvjTVJrjifB+UQ0AfZOEx4uom9zPHLL75KiYmbccPUAi
YqcSDICuximb40o7gxhl8W5PZBNLXbSMGFFgoRqYSFqsNx05LPMM45vXB3jU8icDc4jxH5hxqBhh
PtCzlFJCp472UxlVTmzWOUKLcRrtnl1A5vsiO5bwVGAF2ZXvaqa7eWQo5Bvyl80l0CxC/PIcNYev
4ByS4F8Xj8f0eLDJy5ROe1sF/WMyF5hTkx+K2PMc6JzICUzQa3irpY+fNjRPVtJc/nNrMbnvoCa1
rqjP+JkWpKT0/RLoNnimxc/1SOQZef4BRFhCGELUZkyTp6PiaIOOXudUGXm3qoJ/0FCXpr2wm83r
X8vWNuqzip4upNMeHoQri8XHu6RyafQEyUqBvJ8OTeFCXspMuR1/H9sOk6FGs6e0H03jGuK2IKm5
CV0VI/B1waX28V5tB5sZEXBoxkOyFKUn1ujnaO/H3ha/HAMHRhZ20Yh1iEtmsRz9a54fo/4V1/if
yg+g+Ywo7K8Qs1kIOQLRyaOly0HoUz26OImh2igmOc82pfvK9ZuTnfeGYDLfCgcFJoOuNB/HtbBo
9wwTyNTBuaV6JyV8WlppH8qtW2bIGsnNPi+1xqvSbHkeuld1M1tZ5xk1u0mKzMh/pVf5EUIemKuy
kc/bSJlrnSm1FVASKMRUdhyIFuxra6uncCqff+JBxJn6+nWPRqQYUsqsrsBwyz4PbbjrSjQ0EJho
0NQgNvpaa6JO/fUhTOLd5Co2YGXdbUEDMi1a1RM74jeU6D4QAc5u3pFD0xrNYkthNYLzt12j5+v7
MXUsu1HKS3qALqgyjC1/tRuV8U4+YiL52nkI6NmI+Q/uBec1CKzKX1S8EbfF1YrlAN0WgeYlGOCU
q/BB1xhB3IXlsJ7iQGF09Lc83Iqewh30R+yN5lpUzCxIrSs8PJUTVJ5wgakMUcBh4QQS7tNe1D5G
a+YmwrFBHOWoAbHClz3HfmVx7CfybGPqIB1GNAoJKENidBAnOU/m8JCRfgZ1QEevVpRzUDxn0FGI
XqX6HMW7RKuW/1m9R42OUqsuJpGmgqM8X/LifNpQl9/490HSn+d/gd5LKEkeD8QiOFwRPpE26h/L
xjsxb9ML7tlFMB+ssk9pTHn8UlAkdmNtRgEEv0ndmVLLavhgbKD6Dx9VnnN4l8q46l8aEEZG+qu0
4/HsQPYKJRTmmsxJHKLmTBVSg8IU7hTg241FdA9XZPMhEbbKUknUaUmv6n997QtJ/htHSjtHd6gZ
rUMNohPUsLbSnME9EtefenhfifNKaqU3rELY28g8C6rwvem70TBDQTHl2/O95krjrOz5JB0FMVBm
LqBrz994PvzaUUwQAx/VWbVylJ/5lMLCQEbeCnBkmIxPXi5SrGpm4Bq0R0XgnWSiBlOQQvW9xdl2
HtTYoBeZvN5W6q1nDfZTDS+CEh1jp00BL8nvP1CdUO8e+wGvZ9l/sDLeoyW5gU9xZiyL2WzIgzi3
yop46+HakfA/5zOmi0j8c4VnWFMg4FMSWRwStnSdn8wcj0EKrrS+UsYXaaJPdSXPEuiKtRcsctAu
6F9wBMrMOsQj+YPyDyM4pQ+Yiffm7pLy+w9HE7ujGpJsHVxH4PFRq7U9LHRNzBSsJESsw3eIpZaD
ZgH3rjgrsYNR53BzD+VKuCAiJV/cUUXnLIFmENTGhnnJiIok8iOvsctR3ElQhsqpuzrUnDRaRkT2
11B1wyIdVkQ+fAot5RIJXRaK9jfPt/JtXRIFQD3rj+TxnbiQAx7dALgOFRLY/Ipim83c1m/WlnvR
3Q1Y9i+gmPa9yVmwAPXf7rdWMP3ZqX5+nN5XW+WwMI3kJx3aOo9CRP4CZG4iLkyHWT5g+KTCtknH
UgfM5dqaNrRMDERqtfuBRQk/P//j4WxtOLHHrmIVXorCU3wPA3NR+ASSFtsToIn31AFIIz/Vpfla
e4iiumHhXtR2g4AjIQUeRB2k4EHbYeqTPaVSKLtaQIk5f0jAM3BGWkGeUMY3Pz4ax5BzxI8eiXYO
G30CRxir50Lyj/UYidtmNEtP0ctb0whKZtP9IDGmgIZuZpQAU0saXBnlJB18fQkGdI8FZfmPoNKa
Ja9gF1EjUIq7tAXAnFlmaNtJwcaEROU+9ZlyMnp3jwBuegEkilNLoSgyRT3qhEYop9vo0EcAhAt/
pLccgzG4qhaU+P+dkzMJ2W3vR7yWG02v8Lh7KeEb/LR8LOy3b+SfWVWeem28sQpTVEXByGOSkLtH
f4G6sE46nG1YClq3JNJalZ3dFqE1dBGACTKyGTptcgA2orKaVZlO09t1dI1a3T63MMjxwO9dJJZ3
rnvEnbmwYmL/hALDXFNsFF8prw0gfNrHIygHFll4KV1U8hmlIb9EmRlyUNbSJG6DBjV7x2kZQCKa
ybcZghzrqBxDXJdVZIiy+AIsdAzUKQwhL72kh0Ck1zTQh0j/9LenQePsK1XylDwskfxFG/py3Er/
dP4J0sxJaXU6lnGfkvoaDjiXwFq1vYF83EYcfcrZKjrKB3eywFgwrS8xPVGyzLyOIHbYpQD3Zgy1
EeDKNQSgaJ/nX1s+79So+6xXe6yTV+JUmcJAoVXD8XoXp4hHN5jf5gn90Fq5svsF4BFHD1kz1w6u
dsHDiIJBHtvUZGMNXngX+SEghJ1K+g7GDp0/sD9jNuOCpdlVAZeyNFsj5j/s4Tz2qTrAkgxi+43z
Gtg3w+NLDpcQXvBd+zo31Wmu2mOh0bhhe8V9el9/xfHF52cVUbLio1b+51cfJC62cNCyaoDCXYHD
m0qFEGZV/QwuNP6ZWkXrXvwf7FGTW5NOxqewVbk15g0wmoVYyo3EEbv7fcpZ+sXW9CXQFB1tutni
tQoVEIdDtP53EcTrTjWPimRuKQorI8LZQ/YtTaGoLcDHLHaGacSHn1xLEo3ehH4/FZvhxUeT+It7
p6ibZXCK9Juj99D2rj9YPXFxoHZ/wYyg06j/yvQtRGwlNS0R3YSzWVMYx+6m+ZWaARPQhS2waUnT
djnYTIwDAyhMIpHH58xsfXCjWnFdjI0rt1VisioHrJ1EZiODNdl+pSYh+C7MuyvS+o/1/bInKJSF
o7dhnhZnHHJXv7v7ekCBTuj8xlGyNguOU7FT21vMVMaL8oZSqtS4Tj/GJXTrjtSxSu5GRlElrtY0
d/Qow6dCGyN2cWdFFNRacXCCiHTv+kQl/wNWDgcwVdAg7SqrR3p8nvUjtMp0RxiqP6o4dzMZAHlW
utcOrEuddfTaHiKew9I8bfoGF+uEtLkbxIDPi+nCTdBGCJb8cmbp8gb5vWJgTqIBuKSi6H9VmKTv
A01LyXjEJrhdBfU+tlhDDb6GWjQn+XvIOe+4RlBY+WJBiB7+CGaGSrTcjw6Mq05u/q2m351f0SF0
u2BUN6Joitx5KqJM//p7qKCTJZsjpM2XXedCiVMKQiFETvEgXVKl3v72Fz5z38q2GhwD/rfIXNst
gQP532KfHXzJEQm7TRZHy/5jtlcQnUGRLKxDLv2oIHjauCzADWZbXfIGEnA9OoDHfChEYY9YjCzl
HbiHCdLfdXelBxuJBTvZfb7vuLFcdGh3uWeIwI4tSSAtx1JxmMsR9MJrwuVQVrPKIkRudyqLgE11
05SithTmdutstcdWA0GEkkxXkrctSsO5uWhApj6ImW1I0T1L2aRi39pylwixGlBizOg2h+UkMJJn
/aXeKNgaNKpG4uM09teNekSr4plddP7rfiwyaQBvn00k3hSqZD0BTsV8lyg6u7z8AXVOnfQ9jxDz
Dgq5AItUXpgvxW6PaYFR4dHv/v8JGWbw8PMw7sL/QSR5AA8aWIcxNjpH1ET4mJRAQivCo5/8aR8A
PcrpM54I8dch1/WAyPW1XluC79OgCl17XPxHVcnVICLz+Gdg1WiHmLqRLncc2ErEuB6UWeOFddl3
ipMbBreGT2FqQ6wVlBWxX0UpL2Z9YfNBjs43CjKfnC9o38PTCerTYXDu+twU53k42zjuwNPhxZIM
F7wp1pS8Yol4MkWHwIqZ6EnYrKZEPLOMGSePzwZoM5/gdAcV/SO/Ng42En5MqY+ranXtdud092P/
9JLdQzFyupttuPkwz65rNzyG4MT/JrhnAAbDg4XIl8H73nOZ+iF+u3z2dliHdHNP5tUD0G0MD/zl
akExx49lN8SZjtQmdh562HeU3veS0oPuD32YKfJQMIwnPs437BCFGN/5MsB1Xu3cu2u5ShInUh8U
iS7vjkG3upluSmCa2ES4aPR+ApFbR5trub90fT6HLKOeJyuvtTa9BQvrOa68GXnhq8vv5BpQ2W7E
rh/D9iQPo/C0bnlMcVjyHABZnqzOURsycO1zJPzr4BkomR4LXlsZIbCtljXo1V5TLjp91nRrR06w
dCAjNgvCxN+dr9SzxzsXyI0D3scdjK50oy4so0SvEh1u/3RqfWZHYkBb8vtOWUKMUFs0nirACJda
6Zqloj9mp9nFi59XjQMELT5fWk9SkdI7VFOLztVOymyx3LQXQ+J82QtJmrw5D7JgZQ5v8iiQYWAH
58TtkCaRfjrAIsGNBMIXprWf/7jlsFuBHSq2LFeO703XJw5fa9nsMYEavnihl3YhvVShRN84VczJ
zh43+Kiw9KRF+lud4sPy+PKHhvwQckUxZt7cK/9MOJsX3iirTFq7akYN+wRygfGtg9zTbBGgqmeo
sQHjRG5h9iycASvgYF+0q44O0IyfXIdmn1/p5nS+hoEJ9og/lIHm4cx5t5xHY5XRXRQVlU3Jat3C
M15I8eGzYoZUAkUUZ6LoiW5f8o0ihJzitewNmfACC1l1kABNLw0yWo1Ba0dz2ehSmVDXGQmrLUzX
HOBE8thQ1bDx/pmWfAlSRNylzt1JNKjp8hcUyfEeBTO1/WY+7rJ838B1GEqUjiVVDGM77AhmXKSE
rH2fDQ79GX0Tyw70jn12FkABwNhlb+LHuA+r907fIB2j68LqSuN4a81Mt+kDxhfsMiZsh2ByZ0F8
2i28aK4p8ytxA3B1jNIIO+tpzY5gz2N4xnnm0FmiwRhLFvH7X6UrQNOjbpaxg52qve60edeI21IP
bnR7lAbIYsGsGy7CJAxjpZsMamL2pGDBH+ZO8wUITW5IWXIf/VOsLJ418e0WcNwEdQJZpnfHnR8F
9ArMElclIDEj5ElFnD5ig6SQ+4mlpph2A8K3aMEMK2phob/STnJzDGktc4jKnjJBEfKrEL5qqitO
hktMebADQrARQo1OSliMkMO6mP9iUZ8RwjZQQUqNxdamteyWJGVkr7Bz3B1mEoCmwunDQrl1JG0z
V/3H2dN1znavMgjz+Ec6XKPpLugJHgYa1RBYPv8Uy+qSFtQ1YwaRy2nLeXi+gX6hn8NTD1Ab/np4
Xm8kIpbPZEgR6m8CuuLea3zew1XPl8wjcpz8SQmTKZN+Idkkwa3edHEee1sXoWsdkST+d7NUVwKi
RC1lpOfzROID8HVCWb8NBoyk7kZhNBVbGl1+Hg3VEoD7CZCVOfHiO9fxTI9X7z701eUveHu4cYBH
00xb5dNrLbF6SnzDi2OzfJia7zQzkKQ6QhbgVyxnZw5WYym1La4d9UMiQ2ARXf0ghJsXY78+lvXH
1ShdRDO6W+tVwbSatz6LHFmxXdOPDutQmt0dhOYr/PpmelGqyLPZ/8fJRYItRE/bWA8aiKZgEdVX
oKO63kfNbcy8+yOFvN1ROA3QmXBBia8/EYXKrFvl0VUTVpHSJnWQNqbCNGY/4hqGXhUmdjLHhxKs
4CCmFG87B96ThJGfWv26hQHhcI/0ijr7CSMWhFG3pZmUEVvFJLGC60tRcceMu7rjHXxAPARvXb4l
coax1PCOq8Bc/8vUuIH22wiWaUa56oqngnFIcLAXGD6uA6fR/HXp36MQQY3DZZICp/jREvwhPO+D
mZda5llZc2hc78j9BFsjxjkNJbKXC8suBDmNvuiE4d7HAd/OPaIUfeBAJTtvAfmDEg23m+JkDaUe
WZ5kf/QxF8H7lFTP0qlTzZPyp8BvRXC6nReFTgp9Lpj/mrSXzI5ZehYW/iqtztPq+iOe3KWnaDWF
fS13WCPCb5/78r4VWCA2Eg71Kiv1sA15igXRZDnrYo9o4cDqLfN+mAhZkCfQX/24jvtl60elAKOo
YXsTYY3p6izcwnKDJFSdQe2rfm6dg2aJwGewjROdeC4YqlJQICetloiB0VtC72wQBC4gzMlapLw4
5Tbc/6FS15kHZ2JJCpSP655SxsRfQzPAqTDVhn4nfj0csOnpXcYLlB5kWnajdhl5LyNsLAPGWRX/
YQ8sEGHRRqsuLufEaa8/w7c41Az3r1yjiuANkLK1RniPnNbEtOuLNVOCrKfq60xhMYQWluD/n6xv
nkD8xteC0RXyZaqawfYXIAgaOq1NPIWIH8se2SWLofewwqIDlHnajQgNWzh2QBRFji85tyjFd21d
lH8AfIMuyUPuSK1cq2IwmLLF0DNL3wTRPy97YDFF9EFWUHDlAOjCPGbhBdafxOwhFomaL9IMVtGd
34CwT/GkleoX9/ywKKb1FFK8OHbqG0Dvqjw7cGoBP2Z5aHtiLrZ5F8O5rBLEwKyMm8NikR0YHS+4
fqMFN5Wtq6OS+tXNlGs4iUzpvPj0L8lVHCgcx/hykvDxTLesJCrl0hGiv18069J7JR31uNMrE9zg
gDZ5L9THaMwaDrIYe1Dhj2SLbzUhqOG6wW/crHjjKGim85B2JvMzOme6zjwe0s+7KBJbFueLknUq
3DTbsYfQM01+B0QyrMUUsUe9y+In9wQoSWbsprfPOdncu9ryOYR62x++DahLJ6gOk2dhdqeyVDRC
Op4ZaBSoP5xgGWdBYLeGHTu2yBa9OqgIOP6beUw6m/enWLapMFZVqoEjagBhgq9N960/9EmILmKU
2FWXnhIsabJLU9H9w6rYO7T4XugQ5KSNo7U2bHI/zqRvVfabUHTvLtn3NNhOY2jDjLTfwsMwujaF
gRMnrl+e11Li4NEsgT9m09UbFDaRDy/ZtOfCHNfKWihCDRyJOU6YWodblwvqEcbU/2v2MRgz78dM
ixg9jaCgfHIufRQqVwblvWe54L5D4VjeJ5Hqb0Rd8DCz3hUSCbokRXm/qHmzyku3YIhhhMyUovk6
Xav3SfxELZ6433rcSnrp73OBItDwPWEHIe57O0xPETLRi0sSXOT3r08vbClL2JcWm8ByPbatBU9a
YkBEV7LfOeDkMOmO2iYFQ2/zR/04aN3unNb7V8R3Tw+L4UkXWMY4vXkmpGvoBGKvCRzUZum2Nc2w
rvO58wIlnu01a/dt5GBy76CL9uzsgd2SK7uj9xi/haZk/4w/y0GUB9gOBCbBns8zbr6Len0GaCFJ
mEvWzF4oGC3tPwfceLoCGM77ijE+53UyCikMgLv+/Lonl1XHR7oGPwCrnRMCxbFBg+V31jj6rfN1
kR0vGWQMv1Bhg3Q/lXM6cOAZvnRY/pQdCkFRV7o7Zu1co1G95D3EuHLITkI1g8T8MpnqzrxxTlbW
a1ur2VKAlIe+yMDPhjO2M2lwSU5DDhvhHskFZ6EjLeWmv/tGgdsnZDXRCJpQjCIaDT2LoiQ1SSLR
HHBBuy5SB1O0k4B/htzBQgLyb5Jewiu3rv+pWDTNwQDvY37zXo/XC7ViPsndUECeqFK9xTqeSUhc
yLolGSqlRytecgXPj6qvL/RojPOO17smy/BXvT8jmeNorqgYiJYYOC74lIE8lInXEInKyqUcVxqJ
lbDp/L4joyr06RjmfRiOzyOVM/g4qdAwf/yKRS8sjO0y0peSro9//oQspglAwgAs6mS/Ap/hcfLM
2JQykz93YPsILM0oI6yLJLvSFZIdDVFoI1yJiyRL6hwC65+NGDSxGl0SN8sFW5aa0BYwhyvy64fr
bbZq273usL75PzgoxUJOX114MioPsKf6QdNed/x+6lUzdOJou9lVtL6hRCYb8gcU6xBh9CvXiC63
ivkniBiEhefJgNefvkUQgWK7ItL5KcNyIIUpmlahyjb44cf0MioDWy+5MA8Ni8f1NGaB9MkmXCxG
8O+j9ydOTIlvZm7sGAl8/9dqGMl/rppTV4FHJ8Eie3bJGRn2TD4EGxaEm650IlWbSWTe2rwUALxJ
ir1wPsKHuEKOgCHf8lPIlG9H9RUpNkcJYCR59RIEPTLHKRqvkT62xvnNq7R6GrBVCV3kTbd2AuCj
XgRvhg3RD+Xc4EVw6gveklvSp0AMt7QiPxa5d6STLbMEplPKt27CuW4XAwuUc8a/u1tWzJrx6o3J
0stgWg5Vf6glq0MkTxqvXoe4JPgjXjfpJiSEo2BF4uNafyi94rSLU11gQS6hsck+aIlFpAMDbvzd
xVfHeQXIgkmaZIo4lFeCyvbEEpPsXjPHvrmT7CwphTCuhwzAMU7R7LwpK5J4Mhg/MV5c2gHAVpT/
DvBFJxvVcciHavrLboNLXZZbQ3Ldye3pLLKSnpL64/hJL2Y14OcdypEzfXwdsY+TWXM4BqmkWJ9o
w6PgKsl6N0xNGwEbxLJulnGfLJ+3xsswtRN0f/r2pruOW+z1oClMiEjWufFVscNbVu8NG1KnYAwR
BtIgdVlm9aAp6gxF4cXjI1YZS/88ED+PqLuqkWsNqsE40RL/NeYxNSEiEmDU0b81itX3d6E2iVmP
WAwn/g0jGGriPijIDmYk8IqPmisUIMjdmaWTBD0Xpxs6vTEzTYKLqF1VoTFgOgxYXW/dSMJD2fXI
cGNWIZJaKbxvQQlcXnjvXSC4LWZQIfHTuSmCAjd5FQl7oqqUnUpU8o4Ur7B9k1UisayaKUzV/y+z
99Y+obI//+2iKjCVwDB1HuMNjktw8SJ5jxVnJ+eJojS/KlLyZZeRkExExuacRcKI+wA944iLvs58
xFuNXIm3m1cZgnMzBM2Z2dQ4V1D5O7HOjQ6rphVPKbj4g7O1iyH6Z685m8tFa+cX71QVQiRxoSgO
Y91E33EloHJ/sWC4ThJ9QEuc5wGniMBtlnC+KslT6mVtpo+pTeV/Wq40XfYRKiEkFaUmsSrh/Bfd
5nNxeMKe09bhl/2abgsZo3IP9+xPCimo4HqvxPH79RYkmGwI2+I5mVwzFdJOfpnqNGb2CyFMkKE1
xLqubInlaaakqqzTKXITGu7aKrl6GgjGvKNq8qWMF40T14Qal6cNNmH/PmkrKt+yBipXyOy9VoUa
Sd62qB7Rvh0pOyxpX7bmkEJWhTASs/DQkwAOOr9sUuvdhHCtHCieGfqEwSzcT+pzLOo9f3YNuuke
K9TCQnNFuHz04KphoFFhckXLlnRb7gKMP4YFyEtqAifRxusasTx6dGhx115vZxgoZAEO3sQ9E6gi
5961Lw6PqQ3vell0qMrDmacBIVvGKvydBmtpxZLrvWgc1zuNq2Pk+UcECxMEcQnqndKh7x1kVShO
U3KUSJJ3Tl/d0U3LgcWyttMhxdBxVSQ9sKTrmHffPm33isgeyhpVWGrFGChus/JdAb4bB4HamwCV
T3edDZm+xYl0aebCWneqvUwsLukTHac3lHQaXxLPUcwolH2wlTvmRMnn1IbtYVPAcSsA3wttgBKk
ap3L2nfzqq7upHSKzO5smv1FVOQVY92ER+wG8WBxmdNiWjNg0uJ+6wa685FRKByb9wvuUNhZ18l4
YG7HvbYEvVAwl/m7lsQE4gRHjclwB6y6kcUQk8SgmZcOrE6BmynM/XCKcb7iDZQaV9RAtv2EgPnq
c6Fwtw9Guw95YOLtigussJLFRApQJNZaAXOmY6tJUOxAOytOXnGHXhnbOhb0x17iDFSdXFnP+BGK
PTpcdAkcJ1MvyPJrc/MXB8VxCrDmEx3Sbi8RBa1cWZugQup4iNp0BYbzL5oc6FE0Ux+d8tzdg9qp
xhJCgjok6Amr7PX/ncCBRU5cDpSGPqUe1BrYaOFEpqhHl/ea65XMKIwd1pX8j4CP5a8X51ouz/+R
FiJSUcxzT+/EYhgb+IkfQa5B2X3Zxh/SCc9/hT58TDMuBp1jQ4rjJR9tpsdDDyg9dkcu2OgX1Wb2
bZxnwHROkDwk+Ed+7/mJHb+hc7uJLz9YkYLS5FQgPyTq2ymJji4qj4FrXiG7PYmgOFxiuBncwJic
CEj7z/WHKPbILkfBcSH9t5sv1nWa29Cke3chF2X4fbq80zgu7av5ClmqTrS0TlFrmR6TwGmG9KeG
Y/gmZvyJ1BRn+iu485x+aL46a5hz7h4FjCN83YYctGg7gZ0ZV1Hr9hN2iaBPKzh9NpWZf6/kWwGa
CAPcvr5ptfxwzBkL7msUixl+WBFYhqYoC0XwZK70bMCyVqoj+qyxmm8MMNDtjeNa9XYWsU4f89iT
hp50HHwq68/DNwdjSZZRubUfCQXauWcofqk/AavlBbQtXRncka9osxlrgPMsHwx7z6AU/tT9qKdc
bsjMwue9fiIgun7zC4G/LvhNBT3TGUNXjBpdlPK2+Q22mtton5QbzbFMf5Q3kZG1FE4HszYoOi+U
ewb0VpOLsGLNByEXy+hRYaLsVu2hq7zaL9TPsKOrfBbotNt3M8+jUjA8ENd2ujYqaizyHy3Fknvh
zhXBFPGg9F0k95+dQFiPfPn69EfeZ6kIge2s3L3wcQ6mQGO+SkMLdrutSqTE6Lz/gwLRybRuSEn6
EM/wBMcZkS7p9snQhv3AYucCV6rXAcpJNn+EAn5wiPkh/8Th+GbXL2nGiu9hfY5oqMjEjp+mm8VG
WoNWRQUwJ8g2xApmD7xOhuLg9yhZiZF+xEgAyXe8tPzrnpWAJnJoPxkzU0aQSo+T0Gn1+IrVfuFT
zwo33SJPTNQlwepps/uZNDuqGptAKb+JLRVKezAmjWRq9mzHq7akfTStccR4ZOJIYtdyxxeHkg86
rQeHHU8i9C063wkc9m0JxLjYoOCTE4fI6vc0yu1fdDlql/zbRk6Ao8E6z9958XwGCSYjuHSXzTR5
9+XO16pW/QH47HYTuRwloOrvzEMbStSBo53gW4JuOcHrMcYvZ0I6UxLKyB95POznO35QTGo/MiXe
DJgtNdNOgGZ1ClOlXRfx13bMl2mysGc818fvk44GxU6jxpjmigihXKRzmBJiKI1Z69OYgLd548V1
2CK3rlwyUjQgQy92QxRXfoxnL7Wvn6NEVC73ssvt/b3/fd/Dw0GrLOCGyIEFllpKXbF4AcO8TvKg
afIofvRflvBgxcVhGe4/SUTewYFD6/+yxYQQk1018UWp5sa/GdKY08vAlSpolejDaH5LBknOcl3a
WN5qYG1WXV3exl/mEeRbaNkpSDTkHhceEZQ1O00LanDSiA+ejS24ztc/8wPN/rJIGMh14QQ7cj8u
YvR1CMDfHR0X9oEn82b2Pd+/EdqFNoPHosm4sI0whRPron04H/kIc1ZRkI5xpfC8E+5Mxe4ULqwv
786pEDfI5YK9S2/gCWz6QonKWx/7ix0p1k4C53SKbziPTCkj1DgylG6+/7jxGyJnMaZ/FdxlFcKH
XaUsdeuUpYfhmnOCBH3v5stWp+snCjyQE+z0kNWvGUTjBo/4yPHpEybO2QTOxkFipgPrp1j//pnj
oyAcfYOPkND8IznlwBeogKAnt017bALXJ8uLM8r2JV+l0rf9C72XICNJNWnPDO1Iqs8A3dNDJA5c
izHd6xI5SxiXWL8YkEentA19TooT62vcELsB68J4+IFlcAJmQ6og+rS0/LTe+KMEGZezFJ6Gi0L6
OedOwNfM/DPB0U4r1sgI9dtZcLa/GLh8Vs9VUbk+BZdkeH5YnpFFprg7ai2YcbAF9XK9QUJ0w3tC
fL5tYVwgZVyYTsanmiB196NDymrXF9EQ34DatfwcdgoLtLNgUAzkfp6QbCF4hDpz9kMgZDiw6ky0
55qIGni0cjjjvOIbktpNNl9AckFT5AG0jeMusohap6ZspA+2b0AmktnXNGBPJ9tWlPInLvi6hLly
6rEv4JEIVmshcHi7wXZ8rJ2lFHCHtXKQpMEzL5dk0WBKpp5db++UPD1jl2rOZkyjPgYogaie534r
L4H+wILULv5kBRdtI5B079+KLWsVGmMPcPvK2khM/Ep42MzMla1142jHZy45XgdBlhK5J2FyUPFO
Iu7cvubQN99tktuKExDropJX0KvXSF9FM6VkVSrs7x1Q1R2+gyqUSQQXacZyQRsRHkj4fdjGGIuW
Z46kU7iTzOikVgA2nq7Pa4mCfoVKkkLwctIBw4H02CWQJz9Djik/dex2O9VQIyxDZ/NHqAMAjUjp
LDjrNBTXE/p4KG8LDhlwznV4lqh04lfcDrVZjrT689ckAMbFWn0RUX4FI4bnEy25xT2bA494WX+U
hKHDApOP35mvv2KNNTPAc9URDgNcxpSK1aEO3uX8EbFrDQvdESOZIQTrg6NL02gT+SHHehy1LSiF
3S79Py19NPR4oPf0/JrsPrR0JM5620H4fAjVaaS/ghBERZsP4Oojo6N1JeawpE5Fmpe9kHqmdtL2
zHAYfEmgHwWU9rD8P7AUJYj6tHXq8/YayPCCWcAXlI7xnwrNobb+IWVD5eK43C6F1LPTDGf+05ky
vIkpf6WHQPRh8dYqYZge2vxZP4Q6n4UK1suBXPkRIuLREOT/zbwuUA69ibEupibU/3akrJBKNG/c
9qtoz/nHNY6o3pZvE4qxSNM6Qza7P8qhRFSI6Fn3uwTqiiqQlAwV02fDAeVrCH8Z3eaaT5xfaccO
eN7uJR4iS+tUJLwC0fd32HLSvLDXbjDegQDlHaxr8r4svoqxXiACuZqjg1ijgdWAzg3o2uIqg8gw
Y9hDVI7Gk22cV2W9wNQcFeIEXt9EbYGIz21nH6C4PN9GLEu/DFcd90t36zFdiurtwCaSedOhRdV9
6A33wk7DXZ94od8Py9o7cT/5ynf0XT7hj+HD+lTNDWfGxu7lxuihaHFP38mEHNLexPK8SR/voSiE
haJMMgkFLmbut+5Y3WDM7uqpnyQLA1mYm93Hc0CDtm3vk2RiRA0nuDFXeGmxhBB/IxDWc5JKeG9N
rGGsQVxZaOieTZV3LLXvqQNbDuWIB/8C2k3GVVrKYP8jeOjWDJ+Pk2mnRwH6rQ239CnpNo4tiiCU
LLEAdbbBwHACESIxskXM5gerS9hH7aq9US3G8ibqvJbPdiuPYcT5T/jWbwZghs8+TVkfGLDZ9OTU
E3yhWDmDZvQKjh5J6K+G/J0XJcsmYE5ZV/QbWmiP0YM8qwy4qOy7N0acNdceUy+xeZJXJ5BxhH8o
EfuqVF9nwZrkrWbqr4H6u2ki8bG5QFSEWjW7L8vfSXlQehx3WmndUg+PHrLYWLac3wGAOLAqin2Y
NmizfrevpvvFzMdYr5q/Fnn+SzHGNCkAbAV5Y40XdIdJ6lNon9zoi8X0G9hdqoVVy+NW5CnCL6gU
NFXV3K8cNl/HpNEZNEBw/tp8+nBusJlw7V/C0PZfnqjFtuw45IVI1PRf2Q5v6y2OSW0CQbDl22lu
WC7HVGFY2iT4xTrerzgvM21jXn0+ve6x0ajOJbW1J3htCT9Emnd4nDIzG6wTpJMFLfTvX0WVr+ml
3coCma1UFTkhBDM+hU4dncEH1M7fIcFS+M1PCfZVY8Xjx+ldftz27oT3mxxwFHcFATov2HHSrmQA
guFbBjNFWFvaVO2TcpS5rAJPzo+lQIrDiQ5UxZ7Axh+ozmUH3zMTJrtZs9JDe3xV3aozFdoxCN8H
J8HhOSXrej1iD5H+7VA6tNENSyK6Di6B8CHhjcoDVIWIfEou2m6ciXX3RsdtX471Et+oWqDtdcps
t5sx6KLI/P0j0mcezV/GH+mAaPPsL1MFudKOQcC8VK4YxFN1S+vfZSEdEty/hCwwlePLLV/bgqJ6
acj6CcHzVvk/1Vt/4ZTwmJcDL0t0wnYe1oT6yrpTp2WgTqKkbHjRiFvzhhqggIv/LSQPXymoDWPN
JcJS9ptUR5N2Hp9Z4GAtbZyS9LcXvXDbvNmT30tmn2Ss0dqgumys2mpumEOn/W7AJm5pJJvu8XDx
Kf5A6R6H3lVPnC5C5iTZvXYvPvjYuAL59lNcqxpe3plRl+WDiujus/pkE9g8ywm50OGa4myQJAIL
Xn4rqg6qQuh2YQIcRpJoNF/lC9CD+M4Kw9/V5pueojMYYuTt6fB0sE5rzUePVM+QYLL6tvGTaDvj
qQqf3aZlioHv09tyifAuCoeC0sVnZYuNj1ESkAiFFP4mKEYXbniCFOsKAxkcrusN5mg6WbioVSnM
2lMMHOGk/c5MekGsfo0J00iTIyqJfj5wa+msvPOA/XTH6hAjrFr0T0LjWmpYef3WEnNUkO6uIHFt
6dhm5wxwa0BOMjgFv5cAy5eNCwDDRIHQQKZd51kSZsbqrU5ujj/bRWlaB31apbPVtau8dnODn/kz
/oYTA+2WRiF8TPoEVnfSanYZ9kghCVwx9Xa0+fkAX7hiN9TnrzEakVSbROE4h8bEWfDItolDzgnj
9HiuoMSCO3JM+Td7/6eyJHUvBI7VfEI4LSoeiYFJc14DZI4AQjRorhltZSScXDFQvNK0xQuSvI9n
gGBa0eRwps0rpJFKSAKW+IZYA3u5S6/UsG+Ibth+KmtB+qiNO+W/Um2bM+ejDwcH0Zl9BpGGiRik
R0A7Y5pm6yAKPWBRUC9rYeRS2kyknq4QzivQcmRuPf8WbAykMdq3dQnB51gOG5nW9wIvSTwUg1EE
cduf5rHyz6Q/CUJXySN+nSdkEQx3KtRFP4jNXRsXFaptiEOx6dxCUHAvkk18uLnPguq6k2UrzwDi
J1LUthvfVtTXpUhPut/Re0xK52MtccthQThB8sowsBGZsf/62d1VsiuJFU7zVHLcAW7+4DdtVoWN
4ThqzWwWKL0lT5C9vZpcAct1hEQzOaW9z9nWe0hWwqpimiw2uMZsOMDjfN55v7SeXaBpZ3ZephrH
Mt5/5A23xD2LO7cKf5nNVAVTNtlrYrXVPevN4T7bENHo5ef0MJIg3Sxp3rlzA/rGFsXvD1/E8Eeu
EQH4knVF6CNKzRQARln59NQ2BsooeoV54y/CUAAIKkUf4X3SUlX8U2YF9JnV4a8JY+81XgbvjU51
IElPDEyI9yW3hAWtcB9ZcJpC/KK85lRYR2QqNbv6Wzix8tTvsWQeAE6p0PNlr0giB3BmKsfIgVtB
mkOYF/1HTHA/CObo+wzHx/FS81xeblkU11haWbcXpIeyhfpWdDF0ifzlzvgH+OtPG3ol12ZOjeaf
e781sVtUWC26xDduGEjacCoDIgAQUYptAMAcoyy2Mq5IDBDK15iicct38bvkGtvI8ICTePkBHY/d
SofosLD/ZhipBZRqa8JCzSTDzi0kRbwxwGoxiG5NojPX1IJBaRYAPVftWQv2rstq8LDCcJ3lgOn5
od+rE4prBftZTIIfuTZ+JEbtzPslpEZX//XQfGMrCKhAcuOK91XBcReoGdPfhXAarok7ABPwrcSD
0t4Lma8sufaoEmDNJQOaPss1RTEljYS7IoJzFdUHKTK463fRvChoNw3LSVhnNL2iSLdOzPlQGfMG
NM4YLca9CshSQTNxp2717UVTSxViTDgtHbERMOxbekFUYE2Qu4T2hBYCnTZGsisfsrh0q0jZSZk3
DOHKTjO6THl+0z4eb3390R0dEF3ZMKtaHNky4Im8/xqQgWfp+oKvF6joW8VH7/0yuJXuI9N2DMJC
8CKYnuE7HqX4y9hBEPRea9V/+KzDWyg6i0b5DU74aD7VU8A6dDVyUejEs9foOXpnT4tifLAL6qtu
z4jhmveOCK2Chccu1yYywjQskm+8/GRk8iHWF7s8yTDBCLssgrQZ8P24u9Z2JJ8Rm1haC/K/OjPm
5rCJC7Pao0bsTQ82el38z4pre+zh3hQNwOSMaA+uiMDi9EreZxXVCjQbfZXrEFEtWQYp4VRj6q2J
mDXT6PxbM0ziGPRp0YJI2TiS77YWi64uFC6BhBkGLQQHU1oDjb7CLlnPbSRzhdDvckb0ecFdYjFg
XSlNABL3L4NwEExttOz1UQqSRLcpNcZcD1eVFGEuoGm9ZVhk4E2cInbkRU6NjJx1un7cBUZV+h7+
afUuUtNvd6THGvcTKmc2MG/MhFidgJrUaiSiygV2PURNGymaXfUjH38FhKuITa0m+9Vpa9I7ZbkI
/8QNklXDicoKq1EoZGGlNuWOYSBIVlb+uo2AO4B6/ufp59T87JWAZEQgDAqpjUtySAB9M71Xm4jV
l3E98wR6NSydjl9hdcSwWuEq44De4T48LS/M+dLbAJBPOydem0stWZ/XrQECzLS1PCaAkcLcNXKp
ZSvv8u2dFcsnZSm2hwb59nJCGwNA6Fokv+k/8W+6Ylaq5VhT2IPg8unVljA/TmkeHJphorprDIm7
ygafwojo6wLVo4xXwFi/W5WbfXOovzKU1vlfHUXP0tdraOF5gwM059smI5svrUHIYY+IMohfql9r
80QuS0LYvVAbjq8PJnAqf9WaI8MpH6lmosplMWvtNlnnPHg+FYiSZVlNW+EvV5qVY9PkKP4ifhYc
0l0yE2geR1qyT+XDZGR3yVxVls+VfTgiAVzA4mjPWvc169LFynoe4qS15fphe6AVZZK8lN2224XV
9nrtggy49clgg7hw3YOTB4QSj6M5xwVEjqoSp5q9U+E3IXLY+xtagf+RzMRbGYZJD4XIKZD1fs9H
4ARrcZ4oAw4+LrPsxeNKkezEb71vPdwkAcOuE2blxAB3CaGpGIy66M/iPOhxRUs5zroelXK8j8QW
UU/ql1UTSwogI5RXTUuztNeKmwjiseBHK/oKYqo2qz/hi9FQEVUirmeq3W6CpHn2MVYq0em+FQGX
YX+Pl5K4tbpfqwuQ9+n1pR7RyLpFLz16ZYjhwYGG0Coo/D22Liz1WYSuH8dwpjaggQommm+e6wG7
41njrA8Go7laoeQTrLGgnJADmRQHWynJvwtJ4ZL106Uyzpbh3Pcvrwa0ArEutqXm5dJP/rXz7dOZ
L/+aIqa4bOC4ZTuvPdzih+t4Iaa1fsmoOcI2StAz8WiR2Tdo4kn05bsWdT2y+kr5HyIpTFc738GT
v62plwCl2jcvP3cA9Dgqx9gD+pdxnAnPxlXs6dUvK6dQHvuN8vJwf5OHfMS53q1pLZ0Tv3eUP3IR
eK3eN28L2gxLNKc1/iDDiOCQilDR+rML1OgfP3cspx2FmaHA552vnC1pS8NxLuRC3LCkAWe607aR
kccsje60OyT8YI0IjTjJ2dGTldL2W6uVpigpM2s4qTtQHaCaCgSfgxhRTTi+3+weIV5yZELAZium
VJR2be27fCKJMm9z+Y7ph679CjT4ZL0fcB0QAJ/PtYhZBSP1xY29HS179XHGFysqLq9eoc8NCj+F
ij6EcEU08bx2tUST1XaWqzMtWkqD57+KGxUBO+iRGFPopbwYhxmmSolNIZtksDlvf2FBPwEL1Age
m1f7UAzCrkBO2Mu7D6nVkMGLwZjVCNvxuMRqU9wPtGFFxbaalf4LdH887+fSLOkzSx3DnYHNAZC5
Q+8bkZeojJixbCMzWJxzAY+8mwBuBnGCNXYa0NXvqYTdwpM1OI1+FqsxgfRP8GP6Wy6I3LRttoC9
vuK7cEhQFLOLE+lzczTW5NKKB2XgVwiL7vfKWdiEPO+Ej5NiBIHVmGsOfPgmzKN9E9605oO7iLdm
TtxC++Q0C2JcyyW2296nNBMxmLQmAXG5p2HCfMr4yiVgj0uNITG8E4EOUxig/Dd1pPdDzaJjom0K
kK9ClTtfL7i+bMJjHg4FH/V+AnIY2c3+MTXYfobppEhlLOnv9PR6oFnNEHXomRw8HZQE8w0GiKSt
dSTTAxZMINzDtUC88EgbqsLxPOuBVobNQywOdJok5bMTSVNdKdYOBtE1CNhPdjU5bWfqnBpkUbsV
vNTHMzEqj5YWD0vvQN0GVmILInNkeT897vjpRAwWgV8EjnPCoYemzHYopqpgqsvDi2h4dxF6sF1r
xgBoBxOG7iTRLW2enbSVSS+jfhy00ov6jv5fIQQzFvxdlNL4gxwkoF9a3/K5K3uxuO/ixxTk2riQ
8YBq7AeFpWECzXAQgC4s5w5p6W+y4DFmsb6MtT3OMZsBOC63DMwfD/tZB2z4SoqEnp4Kk9dnvpLk
4yYENtDHlSoh3nZssbtYigk94Aw90hwOheYkAsuBdpeheuFPd0oeM/hcbSmkDcBeYSHqAzYupZFz
42lgsmWrxgx32bncJsTEGNhl4u0flhBhrvHYpxqPRTNiGz6txlFSNECA8XvEwXkPd4JKXoWf3bvj
nfaUgq+3JZaQl8gOP99U1i1eZE2ki62Kr+Mo1iRm7gsMBbtDY63TIhXl4XG4rULPcojS1HoMrWL2
VnL9wJV568M+3ccLZ7FeiXhsypGko5SO1ICMN1vkQHN3iLbcb3AXchnWlutfECId4vDLBhlkSYeR
VB/VZpqMQTuobe9jATramU5w6Zmy3ckVOulysD/XM1W+Hm9FzEyJULJ/cT2uRGaDhKP+8mcHNpBm
pkyqfu70E5pYpgLKrApEuRkk1YM5e5pIXHPkee/NGnZypsJJ2yVqG5/t4VpucF0+NQF7lda/1uRd
0FKTiSh6pfs0g2MwgLC5YeER6l6lRfNJDugF7TmfxZPmDRv+KhUObkHGgeGLPr00o3JpR6r3oZ5e
4GiMsWP2f0Y7463GJD+e2+MYZw2w3rYSzCCa9eDrwyG7vesW7Kaj4is+oHPqGOpgCIoRMvhh0xpu
C17dsJRvbjmOEUxJ7qV1KbIZXg+GZCR1FoxLimXOfiC8n1HCYmQzwPPXau1r/dTKS0BZbRO3lWn8
XQIUfBFuQ7+UN/xI2W06yxkGXBHe6QHiyyCQWMWU8qLbgM/sZlNP+LhJkJDTK4xmJMhQIEw5PPaR
ElLYxZUCPYM/GIoRYgGU+Qh9BtAhDjzQgeJ2N1OfZHFKyBl7GUJSHVnXZwrvO06Ry834IkyZUKIU
RZVrJjDolYXh8yUaaPkiaAaOuukWVC3TLW79lV+eN6cnWD4pSnpAudW3BgFbj0LfO6XHPyloXq2R
lXS6iBQ9gChXeWy0cE6DiNndkRIFoLftp1F3KyfZ+t3n5pwqKNy4lkO9Cfdhwg3Q26nelrhGyzZH
M03ki2X4emIPDU7cubKm2uW9D3TOUz5hcd8CMdAfsDia1XYSRq2T9sBhZ3xFZQEeryrg5jp+Tek3
G59BICtoH0bWmENlOUPGJll+GBZGsDYSNxABJhu4LL0FI7Rqa+sKD4/SY3VB1b7SYXBzD8t+vv7p
EQja/4NJf6yvc8f5o/fQXvqpx11TfJvo51AHHSL8cwx8JMuj5cI2IdCb4ObT/oXAaUkBQj8PDDiI
VXbphIyRa/bM3qu+OOtybzPwR6k8/rlbamskTOHBhMIr8lUmerLdQDsG4TxZrJoBsgJsAaK/IelV
oFTaWFpISpR/pgwjl0VrWFWcMlRgu9sN6EArcWDzZ1Ol/hv0yZGG3cGpZg+tz6ALZbKQDN97SONE
/nBhM6Ul5BrHq2Nd7jx031Ws/1bqamQSxpvQPjZrGjP+1skwLv75OLtinZfXqd9qHEArUHE0lWJH
PTbjGWKNvy7Q6OVzI2Bc11W2kHqPdyOoRqvYRABil/Ifk0SmkNhBDPPAqUOM2e3S5QAeyrdZK/BE
h3DchJgiA8f5K3BNyUbdbFcv8Yjk1OJghpkzsmR5O+RTWUZRD8HRozz2VqWMT9ZHN+ncLutNpXVo
FR1lzVwv3oKXfPhzPuYpKIEp8fF8L82bxlclywtnzJ2heaDc/Ff9n2pPji2g9mWkT+YCmDpZ/FNE
IFUIUZi9Kyygn9Le7y2WO7qrdXLASgCuDifq0mmD6Pu85rjM1XkMIE8KMsjdbfLbczlRZ2A9zyXg
KS5Jh/kGYX3cVyfWsqHikqkLz7uAiKrsfYiebR6JWzceRJOWn9CmqSB21x4ZArt2Yo3YRL1DQ5fd
jIt+OW/QTy67NjRs8g1LVhJVBK20M4tjFAIGlwLJPUNFlj5++xgaRyxGZziY5rWtni+vvDtcJq1z
3AA1M2qATw0mS2Kk9olxXuYCSBX4Qmkj9cWpmLfIJqmDKDoHMNWcStjkS6189AWBjZ6rBulvTw1g
iWXRfXnIZ/HeU7wmTL/jzayY0wgAHk0mUUHtfN2ivXItL6JezfuAWWLOoXREi5qw0ItTeQC8grM/
czrIU0sl6LxoNpyB95zHBoeouTw/dQ8VR8C4jUXMQ21fA9pdObwgAUQ7uYLrZdgFU9kVJb+skMRB
fLc5c3pHuLt1XGLSDwr5hQxgPoV/oBmeqVMP5bte+x8Lyapx4BZojvIxTLbmVMJ/xb2CtuTsC8G/
3HBndwd6YOWSJIeGD31+dGgt4IIXcbEc1ekT7cJFz4RpWHIQuAWqliwt53yvUxVP8zwquCs+Cs+2
g27aHT3yviMp2ovaUHpwHMyhfG97P1oD/gWNM8sD8CSYHbrbU4Tq4BgezjGMPi6EWufNxT2UYxsF
s7m59ux+oo1dM/ON/FTW0Pa2edIdm2q6ehhaCFnbaIU+JXHl6EZpqIyBuPbeKDHpga0c9RlDgGXx
NCZVn5F4REy49EB8cbYXza3DRL2PQc/LvRngYtcgLm1ws8VBEpyt/MY6YlR7XZfEwWb4Ed9nDuOv
jwoHIGUIEBMrVuuJDf62ObDrG+ERWlO9hTsRTWoknKXy++Q2RwIXzl0OqN8WBriRQzYLjIwQC+S3
YxucWt5imhlK3ulCaIq0Piu8EibMZcdrR1SUDhG1BckQLqMsQMpxfrbaRrByRCVgoDAc2tkOZwiR
4kXtLEPhpL5cKbOQy3GPkIk/zZmpAKLvemtAS6Z7hNVJ++JaSqPmP9b8iDUHTg3+5VHFqrbjbIG1
F4B+pH+b+0hkNhTQ/9iS/JpqnjUk5MRAcSDnsZNtbiPd5gBqB8RIpB7gtqdF5DR/0YEeq1T+wxyv
iWkP5Mgm+mpbnHD4TlbJYhwTED9/VyB5eto5eumRMrl6pUcTSBrffuViZ9m9QP3ZKpmPEm+nomdL
pS6RthTC00HZlB9wVcHLA1iEzOubxNNsE9sO6A+mqk4pA40YtHC8ZKEM5kq35VAQ4R5NZQZdtKrX
PcVAeoAB6GEQfxQUB2ep+UgrhJO8FdQLDsN5L+rmTJJWFIuD51vA/GDebBJ9qP6ttBzVnMjqWpa/
j2j0qjd2xaQk7gY3w7Lxt18iH9OSqvp89sG3n2+XFN3nQbu7uOE16046MaIWuL5ZMvU8yf/jwb6G
AClqNjUIRe9G4A8uhXagigGZ/Bvycp2vEy6U7qx8wE++5eDNAcPeV3iGgY6Ete3BcnjQ4NmW3stN
gy/Fc4yKzdCRisYMWHagZRZIf7Q6p6mmvsFXAgdpejeLMTLSthJxhYcsbuB7Z0I9oMCpUv4NjAqR
KjEd1wLltT2zLI60Q61nwMhBqmGwgeA20rOF70QYdZV2y3nlbwuN0W/IC+qzn14XhvcVyrlYeDeW
FCsza+lLhFjKCftncvn51szy0zvBMDkTD4RW7VUGu9dtTbMUL05ld0DGn6Rs0+CUeWtflJTN0BFH
aoza1ZU9dmsIYGi2zuYZ1VF7rAmq+BeN7c47fl2Bi/mzLpqEWtPHgC3Hi9Bkw6laAIEFfTOqVmkK
5ehZ57dPIyVIe35aQMJK6kdO9w8pPUaZJbnCC7zZRIfFHBsGzu2SCEXK7a0hwmrhly9QwGAmHI3n
/3USsYX6+hHps87JeCCk6zdc43+WpGZSYQtEaj3uN6VJ9MIqkeqjHGMAnPky7nHR2kDvnyOiZu07
t7XKWAG4YtgBbKhwXGocnjdnf5MKhwZS0p5uAndJooVYMZoZd+PE/x/84QPE/8T55GDJokyQI/AZ
ExP2tgrO3HRsiy0II9OeXJW1R5QiHcR7k/cjdrPBykHrWl0UgokiDESuYdiV+zQl4ju/VvKmBuRK
bPqJJ+C2ZQVoT+36G/t8G6kLnCpDnQHBiifKK4I+7okXTWpHUTqy1VnGMidQ17ZgsHWsr+TV40TW
oVUMHRvWGAioIu5+yHGhTFu0yLoLbLMS2rH0T7X1mhZzvuAGjiXvkmzsB2M5HeW1Mpxfp+N8nAXo
zi9MiEyZZQJiuxU+dqhHaNl4RNxdk+XGLa+R1xAVZGAdQhJnVJ4+wAFpOYlEz5YUful38BCQK/SA
ktvJl5hR51McWgJvjjjYr3JdC6w4fm5XkIQv0+iG4MEkf9XyE7se0O1vIxqft32AneO5mVZALwqu
8JeiIzw68wT8jkxyWtwN2JEpnTiu/G3MhRF0HtCuy0f0r6m8D8GtQFprwNZksuW41lXi3he2C/Rf
OuqRCKmvrH/D4TkDwiTo/iH+fgmwdcKtcHNxDLgnV4s6qdleiDO/8zW1sIZG7LxbBNWYcmXxTDRh
tcFmCZ21n00fO5dAlPI5ojpAkNyxsOtrMk8+Mb3ojXudU63bFXr0kLdW0XHfRAkG0s9/Jz4kN6+D
7Cije+k0wwHqju1qq9hT9XmOnJawCN1aSqSChqFVMfZH+/cvm2aAquPzlnRhMrJhqzRTMLxwcIJJ
xHVcrnbHYKIpw+5h4jRfGL8SP/MenU9cgVbc72akxQke+Dk/jaghCnqVUwH7rlnqhJXw6nnFv4ny
6LAVODEVy2QDskVhpoDT8R+v0dDKfJVpFLBc9ea6rLsda86fyGRJrO0cHTUoKoKie8VjIhhM6EXH
/aykK+8EWWHBkEwfPVGVtUrEo0g5Hpm033seve2sZ4K/+3MtM8gtDL4DJoMDfgvJT2wiwOG4BE3i
cqLA4vwCLhNJGuw7uHEfBFrr1Sg7zejqG3a3dAKORVz2qp7+ozZU6xYM4SfnwQbzWql1Xm94PBuw
9Sv/7VlnrAVx8UnoSsqdqZC67hxjAwrWNOX7EOet1gwhkV2Cs7meOKhx5VwM6kn60DwFYDTkAwyp
CszBsHjVZoHYK1j32jpJ6jOTmRRVsLox5D7NZOvUsSJ3x7uZQ+I1MpomrrJaJrAzr5/g3XvzPyyu
eFU5vaB/BNMLzeMm/1tdibWJ2tAIS8bP9NoMdgDIhj4SOCei8Fc7yw5BudScPG59dB+MLe4W2SXv
V2gdxl2KOPCKwnqxp8a3Swkrped2H5ZGFMJsykHOuhSrM88XWnk/KE4o8kwreVPle0l0lJmWwgrg
4yJifB4qygHSq6vUiQjzNYaG2MgKp967rm4sXWBtNlJ5fepxiKSqcfUB2q0Ld8kzIYNjxc49M9LQ
ppBnCqmPBrLKEW2JcqKHAFsZnUSp92gpODUb6mwrN2avR3vmd+1eBK13CAWAfvoPVIb7DUFhosbt
5VNILofy4KanRv4ZJNU3wIU0H16lZCDJ/Fy3N7cXXBTxrhJq+5iaZSXnbrSHEhY8/jCu3meK5mMz
oNRSFsXB8IqKeuS1WDST+nWJBaVoN7gGAQa74/Z5RPt2n8YQjepeB9HOnpBsTHh20YdknJBN6wqM
JFQFegsxsYeGdMTQZ9jKoYnOXci+3VrvAjHR5pnXktmPK+pRXFKGaXprbp142iYa2XXfPSF2ZCCW
rOM0evsO+1cGBXz1AvEkOJhl1zVw5Gjq3Ji8k5ZcBeHDD60Zk4o/BuM2xvGlFEWCSUsndL2HApGD
YFIL6D1L4S08k7ir+X4GAmNPLcFrr47FOV7mlREngJ3PuEBc7LwL2o6kOF0p/5WQSttrPEilnp8r
+3qVj9oae85NRvaNYvyVEoiwnwKVIumDQALLqA9QuNeGN3zAIaAym8ZmHU51O175f35BHCTwsZlL
Y7E9YvDVg1ArVlPpqctfjce3krgLQGmTh+H9MBtDjhPdy7egGy3ksK5uvNq1m6S94/sjEkpqIgvM
uflyRT69R8UOA0vtDVe9ovnQfioZDP5UqSF+6kJQhUIHmUroXj23bzNubTGkn5eHQYMrqF0PW3XL
OXY1sYbQ94bhtFeoaynTSx7EhFzRSmJp5KY1fzmlzV1xiA38itJQQlIlQGrl54veSl9kj/6rHmrG
3NwSkWGwdaMQ28WgkXZnjhuYG9rr4CXIk65Bdc+mR+imhV3/TrIbjdQh/0tKFkq0fRig4z1CqwxA
Ex37mPz5phCozgr/6ZBry8Mox3V5YMJIUVRdlblL7mvhL0x7O2FVFGG51miYG7kMe3v8LPaclrVz
kbywKmU/j3u+ZJOT5DCYCaD7JO6Y92nUn480zAT+xmvU/RHUXFQr11Yo5SEYAFF7Lrxm6Ib3HK5c
Wq/ACp+0s1GcNOoBVtH772BnEJIIfLpS060Z+vKiFNBzBWW/mTqo5OX+hV+wJ70AaaaCmecxpu3b
/+d4zJYiTplKC1E1o4R4Nu0uVb+u/iU7qHqAY6i0H998gO/pIWZmQBmZ+o8fyJVqCOZTYq5wtT+r
rTryUCuKNHLut3vnPp0LKfQ5rcnUpOrP71Mfuu6uWNOWpBqH8FXZIZwQfuQYmloq73sdYjBVZsIC
kcB9qLlIB/TEMPYoDoNlplLqEW7kZr62m30+tM6EdNARmDL3UnxXwVnej9QzT2G5N7gF2Z+cNMNp
9WkqzV5Mn5wtFso2JIFpOBvWLbHZXNOY8UoIe3oGgjqAKNa854nVj6CW9/m7xuyWT6oxx95BcRNw
lICbSA+yTxigt0rL8uR3rznu8Uz+WuhFS4b/iEf0WG3DLqk7EVvpZi/9X2HdWBezv19LWNxCRNna
RO8FOyo0QuFHwasghvUpBUVWvX/vv0rvO7xzMWCCjTiDvoacFPS8SnMEDg2sVXDz/Wr4ncTO6nv8
em2gT30AFS4RJxHTe0vuYVBNSBU0DGgfogR5sBELqdiQcs312xS6K8/skRpGu75D2bqN17AEMzwg
IxS2ba2QNgzy8OvPJhmwGHe3drakQmIlgF4qEWUH9U1m2jIBnmhCmki9e5dpYf30m2zGjVVSORPd
LsCk+yZkegLgmpr4RAAjgHjl+8dd9IxKO2aYi+wmtZSI2TfENL9BMdGYynwO2HdNNKnmDt7ZKf2P
VbEivf+UnnqH3DiJYi2invf9ZX4m73z3pcEW+a4qC2RAVbGwxZlBEQV1Sga9xj7+5xNBom55h5Np
GT+/Lc20+KpYcZWGvXmYBkSskx0A7Qwk6ATyet5L9w/ngT+PMg3QUvwHfjkvFckCm7VvuHkUuYrw
noOuVC9WmtR0LOXhF3EfGWcoMcKWGrJzSdE0QuCEhnA5V/ywm1hxC5wkKUrOAanX0UwO6+Ounwxi
RkbnT/Car0EaZf4PiPDP0WgtL3xxClcf7kFHJlfaenCr/1tzyXbVPaLqWSaV48wK8f+RRAhBQJJK
Ngg3MwlDCi0nsl0q9tQtEwBfy4F17NhGFzHUwetVBo/kXisxhdGJIO1WHwtE8X6cLXdQOl1iud+A
HkjpnmNbQUeOVrokVFwHOCvTyZ+NTaAio6EmMCD+AmbyTPWjIgQb97CIC7zKPRQAydqEOzqH38cL
ezo/sOiqtCi2+emJGiRc2Ug/wyg2Hd/dul0Ue8UZCULCtRM96aHmPvILEpaDLx8zgUdbjQ+dsuuy
5zzFPQHTjYTw3zojTNZ3aV7R6kgaRUpGDTyZgt7m/TRVMDm0O5bbMgCab92WeE9soPsVh4U0nmLk
l7aIVYl2FS3Wl85V61tmREDGLVaVJcWpv4tce9RBicJpot6MLS4Pd+A26zg1G7wLA3aq2MU1Z1tj
p+Zoz7O8kdjY1GrEO65IVBSMT9OMm0fsK4ulh4m0xXgYx7rReNNSyId94GnOvCUyubY5vzWJkvrZ
Ogd/fC47bzhxFg8hHZQ5ZIhqf3ZV68KxCZWKRYSL+f0DQyOc7WmP0Y4pJTjotdNCjZoOiDqtUcy4
8HU998EwVHwNdXtL8rdZCmOE8+z8oh93yHtl2OTVNYU0KKWUZG6Z/v6q76rZ+cvvF0+kwN9VDVJU
tLI6TjCjwmz+tNxL4JclpICD0NfDKLjBOkwRBwEGicNTs0kiSdVo2ucYtA+souj2Q0q/pFiSzSt7
KrRKVAvf+sp+Bzm1h4mxEAo1eUPrLo2dXsTf+SP4n8lZ24AzVkci+Vzo8HiKbvJbIaPH0RF2fgBn
yOQ0JcsnW91kealKB+jCDhi75J/2ig8ZFMC6xt6PGdm4ZJwcrT/BmvzAImBVZet4+8A1lmeAiTus
gT7mg03WkUcerQebxwvnBSgGqPEzUItRLPRvd8MzxD42iwXB1pNthhSE8GsrMKbae0EH+tT00W4W
c1HVbMR2CNYSYFzS5+sUqGab2uanuLoBtMeB/dH0ZK7A19LEhkt3tpsgOSvXYPChzn5CbeTPEs0X
FkPykPdrvXLi4NmpDrAoC/uJ7FcohNRh7Gi3a46dVcGdFITM0agBNYvgZaHVI1kl0V/iPGhMYenL
ipJevnsrX/FH+Enaky5wc+PgCuk8CgihzVh/zzzdnam5/9qCnI2hpAh6mrs8dGCMX36++/tftq6a
Xx2dQC2lGnAtqWq3r8X5XnjWmMZcrElDj9k+/zZ57WHgu05V9VKHfymHUb1yKG8oJb2xGJAJ8qR7
85KuTXdPiVlpfg9whiQMWvl4ZNBKfZsIEJ3vfFEBtBkJjlbdSLRMkslcZqpLCxNhSfHFuYSG4wfe
Z7KcfOqe2Si1OA2js+KxUJrIg6m+0Vv+1rMJHnRamMzqC/blL4ukh6v79l4b7alRTxn4pBIFto/7
hXZ75m6W/wuBqw0XDnSimYyfpk0H3RTca43i5ddMa4bUHjeugyjPsMYRnj29D5EOgoiyIm91LUo7
zXPhYX3nS69El6d5pu+loSAaTv0xG3cJcx7DaJ1OcXqiKq6zQPwOA0eSmvEaGITIbLV7k9EP9qG2
K/oyVT04L0MpJtHdfPB28SREXChQjMnt66J8aDIGZTVJaXfMnLNE3lgfXFcbFfRFkcIszdlhiAQY
hXbLRyWTsHEEDJypb4H4Kxx1HBgm+qaoJIJx6Hj+Of4iJ5aub/hukDCleE9YKLdMpdCm8Envqboa
VZJxRXn9XuA1E7JNye913KP+tknY2vQUSz8dI/AXFPvzTyaS8xCe4oY2R9v7bFCXdBpmryr6kVq7
1JxhOD27t2euNS4GmhNVFVdf25rhBEMg5GKcPgM/X0yuukE50nYtc6/d2Qf+1qWWI8fuvYmtjQYj
PqT41SenlCD3SXrOwlgjj+2GcW0CQ0dYUqc/bTVUu7rqItkUk3rIQ3wbTKD70UGaIV9GbTZojj+I
Bik3XlLwJO5aqfVGs7/iM17y0AXnBgv/ELsjnTBRBu0DCNC1j4FR6Aw3UHrV5N2iuwTJuBvBQr8r
jcGKoeZlHtmoKrUa1hbXsQ1ydhcyZKtRQCSb+zcM4nvVlVas92U7qqdT9+DkXlHobD6kKr6+zHQl
oPlmYgcnPHmzJwzoBeeb8jQaK2iZX3aJcW4YLAsEimF4kfBmAGQS8ZYPrTDy1cFVe/CnEIcCC3Yk
lZwKbbaGxAoM3FS22WPOuVyovTwm4TjTltHpFDpGPXox8EBDusuhkRYp9y23BteaQ/tG45E1CWmX
mxKL6KLrY3XmEtKDtiLBlYjrHUaX/5HA8ou+lJSBPmFh6NKtcyfr1Me7DHjFIehR2+PGZIiG3mDm
4baxjEYObNwfWSLArd+e+gHNuQQqK4DRSrlCxnShgAPzLvU87j5/vbUACOIoXWOM4bfjUA+8H/5a
moHOB6O3BpKECWhfAVlhlpkQFkT/B9gTda+bf3a4M7RyM6mY33C/NAD7ayowFKylYW9c64l8tRZT
MIIMdiEQKGck1VnylkteAmPWW8MAu3F9Bne+/fMt2Se6QCG78t9S6oiQ9nOaBffdbpmGeZyX0Mvc
k1FVs6VUfgqvO/RLm8bcNiG2P8wshanQ78km42t7WAr/+LQ7g9C7ea2+PeUdNecTty4zffU7XQMF
xbF5T1h4zGQeT0fLVNt4PHEc0PGLhl85yIwFiKfE4ZZur8LuINiC5Z+NKNm5K6u0qgLAe7/rZCve
YZlprgqR0Mnyju//1F+QpA0EngjeqkxZr2lYfi3OuIhULe+9/r+2BLOHZ5cGw9slC9AaH2akpHRo
89xVqtPk1o+FxuBklzNmPXgpGf0/3OdqZczk0S2KTbey1BNbLjxTIC5Cl6LUWiRwe0YkfH1aFvWh
c7OfQnI3BDM8XFzipbSo7+YRg1IdZtFRdM+Iop/5P386o2Q2I3peQyBS44rBZ0lOoieKQfK13tou
E861v3eM3OcRYkeFqUG9Pebhm2y7HiI0Jgd+TM/znEde8eyjsgdEF9ImVM67czwLZjDJhWLID3az
eIhBicUwmzhea+EbBgVMIQDOtmk27kjz3uNbt3YX/xCtg3LXgAxqjPDQWhAFej1D16TDW08cvW7b
lVo+X7jc46Jqa/AuN61grO6euqLtd40T4H0irz6R7WnmaAx/rmeDgF+JZ3TUAZrJm+X4L/SCIkkK
dJyZd1R31MPMRh8VytZlJGNk8wjT6T9juJ1tx7TxrHBoMhzjMNEs0GLiWrqbFtoomTknS2Jrx868
hgx14Yo3CuEv6fbuLL49VWNwsaIcQhIRQ0gULkV6vzLZfktp3BdMN2BARNd2xv0rxaiLL0Mf9mpI
rRg1U21jzOKSVgZKWwhY03dDHM+7to7qtxIVf0qneTEGdEIWhMEwPlzc0BG34DxaTJCJXszPr7FD
ebbvhdC3W8bTHHhPBy3UdulNvggNUmMPV0Ka+nJNdUHPrHBTOoID/iYPO/g+NRMTGDzB3ad/D0//
hkHXj+fTIGdWV9KDMiwvLfZzeqitm6WkkqM1gghonHFkNNkArGegT3MQjGD62ZmjDTGjB4jQVK2s
jCobZ3hqJvMZcG32u8jAWLi7VpNq2fS2DYtOHo2N5vAUuG13RJleuUPJmznQWnqw8IoNREXXj64T
h7s8tvUF4Pmi/9KVD2Akfr3lIJmeQ/0d4rQg3DsEKE+iFw47N9usixvai0EGdrMoswQfnPyiU/jX
l+nyLKZr2I10PrvN7hJ2bDw/IMv8oR1hJo9MqgjILEM718TLKg0ynkrpU8IwalzBy43WxMBMuBZe
pbcR590Okk8L02aFqMB2Zw6jTBxtsH+3t3iI3Ag+C0UVGnJD1MDTc2T4bL8Rn7qAtVoqQ9ThH0fI
dIC607SYkZXuMZHjOUcOWEgsbRg9Yg1R75x2F5Ma5hR1YG+3G18hiySmuvjehPGb56z2AFB+fuEH
dVP31hLXMtSvCkPUhT+QYF2o+64p5uzn66kLi80DdIFfG1CURGT7oWj0YwEmbK/WRzXd06pvncO/
EnOu64T4ewrEefwZRreAHj+GWQLYzQjiopzVGxejleQOMoIqv/qWvc/53AoxQo4bZIAqvCEEuQBR
aLJ9/huOfVqlg5QXREgiTdGVxBFVaBS39p++YuQ2XP1pZcCYg5aRPZRMjr8jPbNwAh5yndyXoNEO
ncpkhu/4ACFP+KufkU6BPwubcm8U2TGlSoKRw2kGWF90b9TArVyGCk/zeeHBBimZx0e/t2JylzhQ
cjoVg696O+tGQdZOSZX2s/aQmo6J//ZgLTV7mh81//YHLfGnnVZgN/WVWVdw+QASy8DwLdJXu4Nd
A3dB2XeoLEd+68+4InrRePSddFA9bCiIAorStRQKctQLa+UKDX45MRCwGzFKYrbGIptiL1Zr671W
wUGdS8ehoeXj8djAXdAZOnr29S0flh8GccN1wxkU+XD6KYPNy2QPrPXJktJF/rGUP3Z0CfNzuVBf
/c8iU4etZIJ7t0WqyktnnqTlQzKQ9aur7j5JSYOr5HBVeCcz14rdrO/Cxlmdi/YfA+oCLcPixrWD
nM82I4DESH5HevyspVNc47hUdI9yq6c3KAIkMJzCQVgGE8GM6rgtTsDd8wH6NwlEz92Yzbh0dlsF
l+uqU0QWAWrg1N6ehl/mTv1pUfjs9dPLU3ZAmWjDa5lMJQmMMdze3eR9f6566SnUavdHGvPiCLmX
GG6vKBWPztr2wFCSyzrf/1fxCCd2E+Bg0TNjBSjY/z4wJTAVwIURsj2n8ulBCHdSAFmL+3dgJip4
qh5ERW96Cr/5yFTjzrHRigC+2OWFyPu3Evu0NacjWcaBvlpIJF826zQvozLTtqSEbYGJoWpEQa1+
PYFETwAZ3/j5R2JcyXHMiWkOHTFL/UMofknaOpFA3zda7Hrv7XozYiJcHYKOJrZ63mkWjxI/wvin
rhsvmInxxW1rXbzUGoPyClP7zSfhQF6AoDXpJ58OKkzK6SOLs0aGWP1a37n2Ndf3DLlujxLVIF5Y
yGs2pkR/hHE6AoeQ28Xk+CKGTwXnwTJSVFZKFmkYRZImTa+Pzddg5Q3po1kc9lSda3FNAtWEqo2X
jkdjyKxIP1ZMmqJW7a7tBW9JEpNWHN7/0tqtkTj1JZDXnmtF01P1KyyO0x3D8kTNOfPS+3ID1Xna
zd65B9IxnD2/+L+evCynw3X0CgTJWHbeH1+HNtO++dBDTbHCKnk1UBmqXf9Nb+7m8w+QohD14RWW
76lPTrdd4tF7GhsgnkrmQfPy1G4H7tIK4PSFf9LSSHJIYvtmGg204RzfvwOmtR0XsVBz7islJMO7
lzYfgmIXeCP65HD/C/nLwswGAjehmSozmw5mm+5AldeXQduT2lE+krQ71W6zOXJOCUyJEfPlD5ge
JGu4UqkvSrULY6ILzT0Bw3o1WQXdzWbuwKdUH+lsSsHSA6erpjgLzp3zAB6/BBQNsXuICa9EIBzz
4n29D+0ejnuCDALdzUdBlcioNgJ2DSwN+lRxcmkGR/Zjl4oScemuSkmko+B2LvM0NKBgS+De+8FO
TtR+Vta2Ju/MWtKw4gPkTTFhkej6Rr1ceOHhcbIb9xxb9SDREqSoVOskgEYBHWr4Pet106F+Dnzc
1dC1KBSks7jq+g13BIHBCztAVmACfUPpGfoPKHhTiIIgMhgDujX0gJWRWh/XidXpFSrsGLo52KdA
Ny+jqpnXJrHxRHgGLpJ4drh2CaVswN0AS/3k35X5xonIYpAKZ9r/VkRz3/z3luMGmDUZA/zViKKW
06o80LmXR6cFnUfzTaYkTtIWis/stD1VdLF72ogEpem1Uh03ydLzRbPrx5K5sxicnmj9rssl5l+C
H1vG3oAW4CKHoV6at6AgRIdMra5ZCilt4E+hNboLdhyJuSw3naNoL0RO8LZM1NU7AsXmWzL5F61m
rfV5uYyHqbygq9El+F5Z2AzPXAw03FE/o5PVRckciQkRW7NPzaQIXFhRbh4mkUxLNNaEpkVOWWbJ
Pp6noiHu/tGONpWLmPod3lj8Yd7a6JAG8TzTOdu9Sr8TBYralTQDVArcz+Tjh89SPl2qEr/5ERtN
zcDy/dGFCs/6JQYpmxSx+xUgqgKSuNDJVmy8H1W833ZmQCiUI//3O8t4WauXEHAICTg4RuRNlRm9
HCSb4Jfax0U6x6hbr1DgMcT8EM4W2HttZO2O1wbgFt1eSbR6QK4eJdDvLQSS8p0mxwWjEBj6k1PM
+/f+Y46HLhB3uJ21mWDkzYGXgxhzDfG5Sn5jSmoVcZH4uWZTnCtiHFrLTJ3hflknoQRgyelIaGXF
Bhpsp5Lmpzst55vrKgGvIyad2Ck2j5TlCCzyyVK3KfTmvswETqryX0AQzzi+9z7N/w6hgM6TgKA9
Ae4slBEa8rBDDlMfDctzNyb2D4rnQeZH+HDEOdwRZ3mrjlYNofEG80Xkj3oCM/UIh77ynBhFMlNX
ShbHR5SFBfdC3aAJa0iyRVxLKbd/uh0ixw6cMmv7HeS2rfLG4f6I8Qee2pmn8h9UPBy00mgA/9uP
S5vBvQ83UlmZtx+lcwLmVO/SKmbBRzOJc3wlrUYHzY+0QxaLemvXEkEWSrAAxEdpgLVTPOt2JNqW
zBE5J1ZcYF2JMyWS15YaiNPQTsseyDP8TARe+yd2xLGreE9h8SewVIbYuFNc4ZGB5YC2l37mBKTH
ZPbedkV8CB/9Oo/UX1zTKyYJKwhhVoDp2sZqkdEe350WA6v9Xjj6uPwX0oNqrigC6SXV6FPxO5Ma
McdtOBZeg+wjWyPjwlVEG/6FtYhJ1PlmW8IcWKKeSfktEOR/OOZ6XvtI4XdnIfI2SjHFNorvZYF1
vOf/dRnde1fl7XOZnD7B1AKTb60pZXNVO4ylf2XouzOccsOKxzJFmn3wI4Wj8e5JNnnsVBQ8Do3w
8XxKNumOC7OageivjIIqrVj7gyfdA6BlqPrKM5GvNjuvLhUDu5uDkWNtP79w4D6F74dVaG1V4i9g
F9cLRtExhKB6rs/QlnRM8rpznQIjSJfaPHHeYu6Wtwvgf7lrwmv0I3oFGWc6cTbZb84jCUDCE6zA
HesEiivEsBEqplRHYotfL+nxO24qdMKryD+/Qq01qfl17PykLgB4wkoLFZW7UR2Z4X2jD+A2e+Bm
T2gQGImZ12Sv9DoQflnwl3c8pTWeG8xfZh5SvF/k91mvKJTBjAecghnsaluPAtjDyQ1S+EQRjTdw
ZFCxfZx3k2fDv+KopWE6MTVa45+j+bCswZIQ4l4aoeVNK079edqIBj2x32XtUgJwsbJJZPCE9Vwi
3yxZh+DhTTgcNZLqpGV4hSMnEvQgXyfosjdaN6SChVDC9tSqCyxzazkwq6EPPKnXn9jDTzmvk8nx
0O1lKQrh1XMeVNX2o27ZlGQ93PW57EqzFU8uUXqYTWPO1D0Ouhe5qRpfZ5Q3nV66J77hP1dIN7ze
SolwR7G3uo60vuDkIeKItg6Yb5IX0xSgq8qXN5WlGPRtlbXyEpxvKxcf7KZt0baZkESEHL9S3IcT
1BmdCFMeaMfvF4S4Bh1mNxPgYJ7BHGWDD7WqeWpgsCDh5k9R6WGEQZPaLqP/PQFBpDOiP89rdfwi
tvCmPRgce5eAXmE0Qpjw6L2TfqPmH7VkomyBQ5/DikYvAeAMb4aRwzz9JivaG4Zqy8Ckjs0geQd9
ODtShLyH9iPnvkgtAhAYQSyjrjcmA9xVOr8g2EqQs3rFIxrbyL1hrJCgS/qwvKwrxT4Mi8AmN8mU
EBU8854fH78+lralpqTxTPAEuICxaU+4IroSGISHp1UJ0FjBqFmQgZ509szcdldmLLMsVPtd5nu3
ZkPXvl3LFYUaLmw8gFc03oM05Jd7o9+TOzpPxbbC9XKm2LBiTlIBGlGE1I+Xykkhijy8aKgChHbz
PyrMrnl7bAgzCWh0FLfUpvsNrALK+VIyBW76mklHP4hHgwdif6gp+jhDYZXNYcB+kymREGlSaG+p
Pdjz32AZcmpZPvRCFm318k+QHafXRrOZ07ve1LmRbpzoD3wjHUjN0Jgpe4IlAfchnySNe6uXCcmV
JEzwMSxaphFM846ptaYOy6Jgkr5+7EqY7aRer6MkX+4Gd2hDzGeXIF7r++lB3W9HrwQSJBlUnd0z
VN9XkUMI4GGRM93kra9QDYsZvi8UC+pvLxMcN/4d4/BIMK9CqtJxvyR7i7FwoqmbipsHxQ6tpiSQ
vxrT3wbY27E+MbqcE67L1E0T9H3Qg7jOYChbFSeUzqKPiOawzI61IWNydw4y6qMfnuQedpO360Td
UU2neyENRyK8umbGWCwNvL/cuNLK50AbbBQ1Jrk9ChqN6rpdqgDqyw0AIWWouVSjr0h5ctCR8Pqy
w4tGKFsEr6aQlmwaT2T9HstBFl/hhhp4TkItnxybhsh9QOELV0rZBUfVLMSocJmgOZO0j1Hu9Wi9
p0nI0KKqMxiE9IscU6Q4l0G/BSVREwmKj2HwQWkBd44wWOd7mcjHaPCSun7SzRdbFgMbcSNzkUCl
gSWVOJMnRGoT+wWaC1msRt5jiHVID/iaGFWoMbXzeSpqLRBLS3jNMwSNshAkQsGNNeDvm8ScdliE
rUwBwO0r6c8BD0+4SQxS54S7R0Zd+G8ltLRJEY2Nz0tAVO3TInWIF8R8csUzqLq00PV/CMU0T94g
eScRg60PLjInJM9gideG8LHwonINkBMTGOs/LlUfUodhCIZVP5pVexry0CnJ+lUdI8iKD6gi33Dp
suxPH6PlWT8QJ5HvIEF/gCgHkNhJZkhLokybqpEoSso8Z8A2PL9dDxXNC7EKzYzQeRnyJ4jbUWjO
7oT995hFrgPzh2MC+OHHGLpBXpp9zWq5eIZMa6FfTpzfDKAyHOH4SicvBpguw296Z6qOP8yyJtUZ
Nq9C5KEZlDsV4vK38jihS9/YBcPH7IyqdhhaGA2o+L2VKrmy3g4SLMWn1ny4zkvixbycWRd7vMx+
Ioi0p1IwsQWIB+52oqnMliWwCbpJmUojJH4RwgSqRP0pUp8zdvZzpLKZ16MF0q+hAq+ZYlVTXxsZ
uELopeSyb+Dxhoqo5l7LlhLhCLBit4bYzLLS5M+poA+Ffy/TtrPm4fseyKVrunnNfPhnaORmDMhB
uGCDlmThwbkBr0gLeUZ31/Y4dsZST8u2F2AvArwRD2tVYwrP2BgI3eWJwa4tbYhFzxNsjPACv3Ul
n2r0o0DFyHeMqDojIglIHwEhWQlTV5SiOEohWBX/TRCJVY6Q96b6h9MWtEGeciaZFUZF2JcM6QnG
x4BKb/GcE13jnl7akrixgQGFiyopHjOfIJbYzXh2s3Fvp9LAKP8SHulQtA7vjd+O8VITnhkvp72n
Z5HQDSOm92nz1lzeUnsZMSldNwgRHw2mS50A2WeTqJC4Hh06N2DMyHRniVPJHLi+2/q9oOCwE7UU
SrnLL49vpFYwo1+z5yg/MT136XN2Go6TtMtBaHO4VDN5IVZsYmpsqsjeEvzoHo4ggJ+LnSIsgPv/
N3GOaS9t0ikgfG2DZNdzq0X56wVqb3Xy514KWdNgblCMVogZ2mcKghhcV5PgS25mrAVDEHkaTPgA
XxCHbR9NiQPAYr5VFYs347k55gXcfbtphie51JjhSHtMfIahfx3GeUN7yfp2x9kKqAtM76aXK3TB
YZERKXLeLO2COI8/OUHNqTSS5/eVKGdWwBayE0tOgPSvJyUYzcVu0rE+9jQlb8iafOqE9ZmqFl7J
CYaJeU5Tdf2cly0NL4gBFVT90f7kuemDU7pongHz3tzeuP9kqMWzglYCi0IlUrLchNEsgz8S8m3S
DrtiGDC/Ci/6u4Mnk0NIRi4cevp04jYlxsaJCGK+32T8ieK8Fg111uqJMfyBr1OmKK7QmdjCTlLH
+CJnfhqKrUK9emCJZm38VTe6Knmh8Dfx3obeYBfUTbn4hM30vYZGqnHgtQr+BkoDY+/eGqDswbzT
g5Cqg5aQEqb7m78FaGZBVD+oid7anf01dL9ww+MrDkOctoNKK9QsDuBEGHXDCneuHUHCqadoVY1l
j/aFCvg/y9A5Id7/w78dF6mydxeN5HVmH6r3AEz4un3WfPWQRx0KKGckUQ+2W5rtUWa2UGJ5kzv2
tkimgx6LRgniP48cfyz8kCOqENRWhO2JiFHi6QfNw0UuPfRyAZH2I8TTiQIRPD3KL62w8FLEtRRg
3nNiSmGD7P82P+lhNXzuqF+dXEc2UOCyvB1Rs4IbUzw2Fc7KqLzaGhCW4sG7uNcfBkeDuNUeF7hW
UXTd3feLtNbScGNkZXor26X8I+zTLwk2XUjMaxW8hWlOPKfqHptdG9jl56Sj6sGXpKl6+dNB8A5+
RsMy7P91XQiAdhP7juj/Y+HOniyXlEZSLHip9L2k8sU00npe3UWY33q/g0ao3aUtR6dBRjiQ9q6u
s+IYgvc9y2B2rpnArhu16417KRxgLilEA+aE/UjBD3vJdMzB36EAncId+H6EE24WpEkndBZ/LejL
uZn2/zgeesLeDuH/o+RC58jDzgxdxJIUaTW7yAuUfT9ZUdt1A+fM6gAHJTH9Q8RIRpScsdB0oBV4
eJG7klQjb+KHw92Mce+GZtKo7VETx5AEgUkGZ4IXXzgGCLkaF/s0d2UAq0rj1jqtE75ptRL2AHwj
lVYkgrMUSUKCZR3ZxcniPUz31lrq8auTegeJqzr862iUH/9mNpDLffV8rUWFi2XXvk76fFqmyAE8
SSw32S+3O0Pd9aU5AHRXufUa22uOuqrf5xsZnNANo6jxN8/UephpPY6KYJeDT/MJ9Ryvz256+OGr
oE/hyQIEZpVYXNHVBEu/815X+s5YADEMCB78sw1O5DDUBXZ5pPI/OtSWl2GA0JoNGeIS5Ei0jRZX
JMHrDGHaxkzWV6lzomRGJBQRADRcB55pykYqIJowGig2dswnEP6mJQK+QOS6GK0n4iKKGQoIKVZx
XHXZUlDs2p1/nXG1hURIjn98bBmN5feJdOuRGoA7mki8XNJNajd4wjLqHZeVvNuQ0SaRbVFuA8bX
jX+j1uEJ/IjsO6/prWI6zzlFqIleXL3Kh81IxLcjAdqD5X00IGxrrUyS1kFPW+tH83yoho24NcZV
g39nnjzloBXQRFUBHqfBCVNNraLvmXp4srMc0RtdXaRxRJ4opK5qrNBj9xxQfNfYxA0yPLLUbnVv
AUL18E3OH9G20Z5x91iGQApJJYc8rqRqtM9dE1ckGWeQ/QZtFWB8sLJxv76IeHRb8jaFH2kz5/jJ
F6lTay6xzc2O6Mc1NVLjNCpWZ3foJ+kX3jqd/aTl1Me2MJY2Vaj2VS566SpVsp3Ol2Xx6vgqRaw6
/POXKa+svyKKLTdaGWF3eSOVxlmbGAFKtqhbS+SGAYGcWqC6t/xQk31/yronDCPy1bPWpj0lCOh8
KN2jcyMNeoF0XiNBMWfcscEJ27BSJeQHBrSgJBicMb0Lor/6xC3dItSWPWVlPSsUZwb6vcgkCOVC
4G2PODsgkyrveGgBMfevrgE2xDRAyCi6hAC0Cp0Oq6z1l6i84qbICNR98Gi90hGHu+p9uzlzKV3I
DkzULqYHOaliw0gzBFUuWouZ3wRFkxf/slT1M+VtYUP8ZLsPsmQ0t1DOgW04DdxvBpKi5UKmRjRf
QzTK/djGC7mvGvXA9h/Xgq4mFhRgtxi/+RlbpKD93/Qq/bunnipj8vW66seQLkuLSbRkc4oEQIkL
W60ICQOcuz6jXkA0n/BLHa2JgIl2mJEiLLE/ShaQHkS8ZIBJp2Wyhf67rRSitmX40Q92GSfqyr2s
YlotH/4DXUf6X+f6ABYHcVNVtHd3Rh1e6tbXW0UMNscOjQ4e73xeaDVSxrVHEr9sQyWEM9odBBqW
QXtcY4Fjw5gs34GazAivn80uvUpqtEf+ng1XGmpKtUgNtWiKB+cLGVSHtRlYcf6TAsxMBYLTT7qT
K2Vp/v2BXHvfmdV2K/1rRVd15iwO68VDPrnjauxbtUqKOO/1b/6d8tVOh89qOo3uuhZRixfcmmiw
2sUDC+Mhmus6kSxLCise1DNWtHr0QkX4jru7OY/aav3v7lXCh1r2E6iyICS+4KNmxNNn8h4zdt6s
WsR1+OwWN7OYVBwsMqU5z3QkNFsA1yt1azadcqQRJCcJi9taq+tmH0ZQLg8c6IMKDe+pR/uWpe+Z
6CoHfaRmGyYw6mzgrG6uK++08itvnA7lRqnEjQZ/spFb8HBajm9GFQFAO56gdoCfW2OMt0Ayvum6
f5ead7yI4U3DboiPc2rH8oZwr269DpEi5ukR7a8FXnDsUbtpbO88zZ0cD6E676hfq03zRHllMG83
0Y/EsbDpSeHBRkxU/0i8Pk/m521z/IQkMrpmBHILsjNLXrtZwe32T0M6By1dNF4SmFSSS6Dqvfjn
GDfum+LzFUE5vMK2auo7KcbOMCXg/NJBDxJa6BIocX1WNHOJa9xXxyjR+DbMVpAQmz+4AdDSUKgw
0e0IwSzMGSoz/0DM1xvhlajPmge6eUvOkvraITdHkntPbl/8/Y/Jxins0wSQXWTX0RTvHCljmQFO
R0yKqqVn5zSKuGP3cCJ9PogmlCmbmosVgoSzrHeFlBn9Hh3Tm1xC8evRL3YzEjgNUV8Xptw84MEw
jN+Dk2VGZpgYfrNmpA9GEU5h95ZUa1fNme5ao84hiIN9UN5cMclwDwg8NP5Um1IAhpgpQmbFSwgi
KS++KCi275pNOulvrXlGb6pYHLb3DyJ1dZXlpwuEbgHFoSJsqDAW9Cjp6vROvdDBg1VyHcAMbhIT
kzaDI+XvkWAWFanSH8eoLzGGmZpaILLBep/8PCuDXsLs32QYthS3TkkKKVWR+7OlxcrF18ALiPhU
iMAWeSbUa77qGKYQLxu+6fTlTEoGVknz5GnsJhiqvOVQRCKOThsyF4/uj4MjvWZcuL8EpThXDWPj
VB5oAnXRqH79lBwjlZIIeS6rtB/9uUysOLOo+lCuRTYeix74PJoxcL0Lj+dFmj8lO5JTqRffJmcK
Bzch3/RtYoA59JkAY7N+wStpDYbmvidTWc3UOXKnGrXqPshE8+n87GC8hBe7aeIl8HhdDLah7F6B
r9pL0x/j3oBKseHdLH7/6ibceEXhHUGkliu8oCMzCd+K+l+Gt1n5ZpWWgS3qddgDb8SPAwDR016E
nWUnXXevwHixoeXlYbJ7AoqzBYYjk4xu9nsI3ClkfrVxpG2bFgsq+t/UNVagZTR0AxGLmxLF6iFf
Phb5fcagR27Y30Qn2xwLMJndPWLvixhK+/0+kssp8oezZGAHlYMS3l1COYayKRFiRGWzXiEWI8Y1
CpiR4/iUX0nv2FhBEQ7xdDAp/KpEKZ4ld5+qz4lMbGjPBzarphZNFkOECOd6Z2Qz1UeQtT9xG65e
qs1ZoPH02g22WBpYfYMZD/brQ04O1BFqgco84gvehqOYJZMN+adZtgi0gV4KRPtuRPE4YcEUH4Hf
SUM+0S/7iy2B+brOTK0BHcBebWwOia0rGnIOTUMKlT5+SqZCnIhn+Ryv6eiPuvcd27XRWAxjausL
k/E6Mt+0ixHLFZT6IpoiwYMexlzYHRY6XMqunQfcdjnAXp8bBPK9MVvf1XY8HyBOxNFBRVvIMCD8
YiJkm85bSWdT2q+P6/WUR4TErEngai5xcQ5wssd4bjofpSD46IxmTJzpjZUg4qLM8nrxIx63DS+S
qSvaVz7lrnyDcDohXppyxZJYfRyKqMwmWN+BLgxxGmT8+1FWTxCUEmRoiv4TZFZzrgDo6O//2aDz
gfJxgVNUzJe6Ure7a2lMq8m9BeDXvAYzqTbdFOAMFjf9sUWmPXhLzT9CVXy7tVnoYcFzJYDLZlh9
AfqPdIdOe0JC5b0iUn3ieLG+bxcUVkpx5mv/EFBaCFf0zqO2QJnmMX0v7/cGnXC32vVwpTu7uSBQ
JR+W1Pp8O5QagmK/Yn41U2NMx/ImDiJt63ShzQDS1tnpm+8v2OdtWCvjiWzCvO/4oKpYOq3CEo6q
+bFJub/c7g7hO6YvWnl43wep7MBdn98c3O39rbfodwT2jVfUgUbLcNZ8FMgjUYTae2UdxwV5Eo4R
zGgWoMtaLQliEe0oOARnPfTdE7QTw2JPMyJFf3Z2QdtR5KEvdtYzp6htleVqkoWH2Elh7Cab9wSR
Zr+mLJtCCYv/To9hOz/zXBervxfslmtCNJUZyc8a4w3gaXVrdkWRPFOJ/5quYBpNhZ5B8QVnM4Kg
PouZNUGf1HLP2s3cHuCJd8NbMXVok8kUlvlKT+VjfjlpoI8HJ/NGQNgikSuM0whHLzQSMbsZ1VRu
KR4FGgyoD0EhTxGgeoTsXd0xtLB8xZtPu71JD2yH2uY2yJF1tgIl5BZDEYfAk0vyi1rCeAF3X/3y
SK2k6XtIeD6xAqLwYlZeSHRJgrvaMKabE32RdlBk3jdk5mnOD9xBgoj1j9Ow+jO9WsCZZzR5HpT4
Ewjg1VH6o0Bi/FtKYaJfCApGYgY1MQfZ+w9prejvIdnIpGE2BS3i6l9moj79i74frx6qk9IzLgap
OKn3t3TIF6+t0Nu78aCQvgeQzYIDCK3pPyGCEhkuQhRQ32SNKZxd8cEQ6vNPaLt0Er8/XGwhZGGb
ntoVbQFJXwoVVOlB3fP7JdnytEpJz9dMUw1hQPQSt+UT1mQukVr6yGXD9SvpxHXBY946BPy2clfn
BDds5VlZx32T5/7GSzkwsv8f/i/jGniR+iWhRcRezaICKzRA0C0aKKvajdNRk+5Dju2abHcg+j6r
3gylIeWHYFxIUEHX61PRADgdczecfPuNaKZr61mDqfTRo8NSEp4jtzzXE0ybN9OgFjBIuDqDpxpy
M6hPW4ShaNYboqicYep64rREP2qSwl7NLhMSma/zBEQ763Hd85hN1ozwOWuisH3WguFaOr1m8tfl
LaQS0NTbJq8dmrCq4bkHFTid6j116Dv2SWWXayiCDuwBCTzh2WjEs+Rnltu5KX9SfHV9gO0kGohR
3uo/2LU1oE6X2l5zLQNIq5BHObXzdinfvW9yT1SeixOiNsAzTwUbTFQeFY8Bb8CvVXUm5s1/n0Ki
U1p52S2SvAB0H8G9t8qfl3eSU7YFU0eeS8yzQzsYPQ1MSYKqkfhER8i7ts7a0iQcxkliZ9NDDiIS
XdQmL8lkpMY5UKF+0/9jot+JrI5DZA0AnGkr/0xrCMOXMggGlyx5iipj6VlY6Ii9x8a6qAMeuNm3
e2em8DrHCPhOu0lrrO1BGgwzwpYut4suxHIj+5N5D8XwMiyU2ct2+HwV8aqEwYs+NhXU6o3WzH+u
MNURli8nRxvFy6tM591uE9hefEJMi5lSm0dmm4P891snIg7NC9aDFfLdc8qopjb8SvR1QM1u5ptZ
LSoJXpo3S3GfyG2rIxm9afOgqp+uOX8VzNKlXTj21d+g61+Fn70x23GM1YpU9WQa7jKRyamOu60b
GKycj648rXwa5WLqKMtpRZSed6iKQJP+2ZDHtpbhhhB1A4EHkstxgDPB09iEIZYstVpjyl0bjMt/
1hdPVO6YeOCVfSqhycVSjUrgG/H5jFXVt/yTi/astwJMxwcmbwghNS2o2Qv+b4x/5LEQ76DETdVt
DslFiPWhD/UUVbO0mHlwVMA/tQ9GLWvXzmZtFwk8PQihYzBFJS/kdDi9pMzoOvbf6vY+1WJYhRGP
feioKUabKsxWhvUJ9WRnTI3ITYxL2eo9q9ppCkpj0WDNDCLdzK9Tcx6lYasBdMg63ETzmBCYIt30
7iZrn3PRGIoacWIzXDhkY6ewg24gYYY6bQR3+vzxvkjteyek0IGG/NFoG3e3A4o9HYuOyr2yktFp
+kykrv0WU/03w99dX7Ym/Z87q5fmuOXIHD2ZeTbDvobdfgwuoR4wj/w40ARqGvBNRATke5Ljupoq
zn3j9/A5Ym/u+fPq39gGDouwMuRsnz3ga7VWG5sdLquXbmjdSSQsHYNjzkar0yLCNHyiCmnUNd5E
Jer7ZiqsX86oqsH8vTshYZ++mD5kHfxFyVWwPogqhFuKK+xIAw/bMJ0FuZPUIWhoNaZkO7VqUkaB
mEfwND5qn5F9X2i7dibtmZDm5/f0vKY5az3eXDY1pPSm5Myf/cWe1a8ylaOQ53HBCbffHF/Ygmig
gagc80UJdvGzk+MOwd5Y13vW4wyKJaKpMRGtEWsbDrASi57XGb/FuqVT6STMMjVwMpIeiNvvfYUt
J2JAs2vU6APkEWuL3WxaHH8T+T6b3QregV3DuAhKjjmvbpjJRyqb7HdgAH1I0MkWPws5u/hPzP0V
wqUtGo9UjXylpsPqf/mMb1gEN6wPWaeebRBj8X72AbdSSrCQ2NjbRouNiLymPAOpilQCUDP63q2s
Xf9OFjAI0dz+36i2Yh9yPfYw0gXIIRfmvBwEkeBf6D+KKHkN72jT+FdDbqhzdu4kNxQuWmuzRZdc
tfP6CNBzmKA584LtnPrqV73HEDshn6UTEBtkTOLBPnfFok5XV8q3nxSi2iOJxiZ2IX4Ev6FDGmfe
aKW4qyrwUygqYHKeC4/eGP56ZwtZxFn/DR0Nr+RWytpDoXyrFoNpogUHOU5iE8nTa4rQZm1lXMF5
HFwuLWcV1RFdpekS9rGNawRMfNjWTFje3Xh+o2KZDsqJgnAEA/Wby7UJomYS+D36SyNqDa+8moki
hxGMQMG3Dzwy5Wmteky//auoXwY70+aPjYAILSNOaFoa6p0WSOZy5c1b/WMj14dvvgHD5fnkETfu
R99wDtaB2m+FbLb9iPTT4C/YzRNamX9KWEGNSq0e3ZICCJHeXFzlLOCNt1Q858OB48i5Jbj8UJdE
Xe7H3u+rXTivHmPUfe+7f4XukClbfIZt1POiOGtQT5iBbT5WNYUI/VHJbLONSyXp3NdIax4hBTNC
QUzVwGaJ4s83f8qaoRRE8KGM0qFK/sXlE+pTjCvxoNBw9G7MaUSEDJPQKQo1sqgiE3OlaXUFl2Bo
AfopyD+2u2kog9PXQWJbIwXPXRlOIuWHIIF35wtjRXfuL3SQKmU1YW0OuZtvu86QYcpOIhfhm8Rf
862D07k9QP/9+sanVYjoff3wBdQFW0Okk6dy/gwiZ9TCpWZOToLsNZ97/BPqSdtHqpvh7c0SXq0z
afjzGwKCYlPf7J2QKV8ypN0h7m98pTAIOBNnM83PsQKKINOzHC6AkCMiKeCUYow5yfu1XW8YXqWT
gd/jWzub3fU7FFIi/6Nv/CK1BpMey+D3kTXBcD7ImHhdd0ZnQYOk1VTDBzD2sEYyjRiJ6PQuT2Yz
V2EU2B76A+LkZnbfcHJExZkNufD16fEpELswe/6feUbakjyVHWhdxlfYrksxPINRq/0EuG7/AgO4
EkILY9zpc5niuvFX98g9d8ANjqWrX7FxeNGJzHmkfchdNruJa6HnOMKBXTQxL251Fmy8m7Pou5Ny
Z75CCBwnvqLUDfRHA3j3vZmD5KvgKwNnEwa4xmFe5RHto5HvJ0CM35ogH1rIa+eSp7FPvKnUE2st
6zVxt50vOnTYoaJ8wmnAYqvHVuWneMslqIJ0QvFbVfeLAcbHoGS/1NPYpmRgeRvh9A+HWpY0wRGy
h+Leujg3uaszNxROwol/byEcYbjCSYusQ8lKb7P9/IzCXS+1iYlaEoS66q14dBIKjjDB+p+uwd4W
H3N5vbGI1fFTdKpBOi5n3ZnX9u1Iyf3/3dW0oNCcCeh5yYsuzqowg+lcut8CSDyu+PxgdEgEvpTs
41h59oqSCkUpL0aznNfeAIv4SsNkuXGXFNEblSfbdSJMVtqyDOYx1qg0FHw9PGRXGlJGetx8FILT
CquIbvfR+CH7ZeCefGncQt9tDwNQP1siRC7BbCmnnmdOauNhy7nedYQZBTV+EN/G+U4G5MCmEH7/
n8F6UPnD468Wo83Q9eyfMwru/fHX5QnxXxmgm8sId9G/m8Lc2VQI6ImWEdCDklffXKZfL/nsidAg
cBiZyyB7X0tnBoiOn7KDx5wcWifq4kCnCcbQZqkAegQT4R0wfDhIAZDaIugyJl/CVVqN227iEkOW
sNzwYspJHQBNn71jDp/IU9I74GkoEwozlm1zENcyImBow9FvBqUIx+jFVQRVHKQr12p4qtE9mXjk
eJ5e+LETjdQdkTlBPNG7vXu64s8Yb9541AI9br8Iw8Q1EfrE4mVb5LuBKBupGplq8BoOShbwhrum
DryB9J750bPVG0YjmSOtCfR/hCDWx8CXLIvX8opttWiQIPj7nhX1nt4qgh84yLixMacG4ovADMcO
k8TpQZRlDt9s2YJCsZqaAVrvbelYdo/YIu5KamYj+AVbWW8ndGd+1BMi6EQQO4gwjAxk6EaeftfM
sfatrSx2I9NlJ1Fd/YsSMJF3LRV6TIPWn9FoRtEZ3BEj+O0vQaD/R+8V+ocTvVHtYkITOzQSpXvu
lJ6ww9MS8EPZo1tcb4A1jNxZWcHAoPE2pHciStTI3XKc/7TJG+C+VM9+OImxTbHetgc3ehI1Us9J
YPQdgFfmRdjeskA2KMgGJfK28VjEdou1w+sv9cuWecGKMdFxphRSMlvFZ1Sbw9T/rvG3GLyE+Bwc
vvZ7TlX4l2tqTyeHHJX9MoX3yrSqLHmxQw1YlrIzvagaychnTS8gMIE0DTdWxc1boQcFbl4wLv2u
fCoG5uNCx+ISakWPMvBP0/CBvPwgAuTFcpS001gxfefWKPKwHlpFf4xk1ZwYICA/UZ3RLMqnHMhU
eMsRI99B+1YNGwcex7OaCn3CU1LVEQcR7yL/n//tG4O0EPRAtV6WKQCosYaGRMCyDWNOW8WYh++X
6Ow8GBxCTO8U6EFXRpdORwVYrCsN9kXJPPnw9PaR/ocPpxr3tgb5/R4MoepHZmwPYLNYW0/g0p1H
Ws38vify6k6lekoU82+6IfGLBBjX/Wl4hvoZ++xGfEC0EMTfvb1wBT0DRCOqCToEpml3Zrl1rSAU
ByTeGiarmjOUCkwZKcZFOaZ+FU/kv2e9VwDOb+GYe1Q2KpYYT4VI9tXTKhN3qzKkNISTTkUnkvz4
oyRQGJSSeyWdtKUsqCdFNi06nWeasTO1dPSmNbLMgwxapVeCQuCJwTQZUBU8TA6psbfvWWXFYSJd
8Jz92nlFwbUOlhjRNjO/VlPA5D83hISBirB9hytNSf/nvAFT5G8BfiwjplFYqsdG9qNrvx4HCvVP
/dP4pskZ0C/0tKFg9jGMAstbK2RRPQhUxgQwE7rZjWuaLUbb8hoE39RGmjEpaWUXik25zK8P1liJ
MMdLfrKRr40SGxjjKw75gvvM28uEDAWS/7dl5rUYf5p5zhumAEB1yD8j7f9ySx/lOVCUEk8rCwtZ
NENctg/dSKilyJ443mxiuMcOQ/goCXSeyKMh5PTNZY+OHhKRvrjNZC8U8cGW54D7nXCO3JIJ1n1+
1ALNB34hMDX2nT0bkEplpdFNh5ji5vLyhXCmN2vrPZPensVJWG7+PKB8yHEPqMfhWCEUc3Ds3+FP
niNlLZ3xPWu4qTFSvTuZf3YKpqVM189Ht+7q0sjzp9pdfbaKCdSdobPm3xBg4x1n9toHruI2pcts
CkylSEmS+LogZ9lMJLm+gGNDuZoePfSvK4NQfO0ln9++tqeZKx1s00kwWZKGkJXVLY2p3BLKu1Su
Aq9OdFO0Drxf3zMtm4luL2tjBwko2GR+D6kulE5LLjc1Tpvy6oDE+nwnHPIvHxJSVLO/1BR4Xmsr
4veR9aiEF34KsavY5KnLN/g1jZQgF/gsumzxr9NCz1VQ/UdxiGhwmMHROpAdIKWRYACV9lxxAsok
YsmRXdB6laKyGhGLg4QWwtlM/5phvAlI2MPenwWwlRtnMMSRJ2cCrp6YVU8/Orbtz0oroFNkLCWc
cUE6/LgPrPBmSdjpOPMAu0WeSTpEFS2J5GZXWccljv7/pPmVZ9vJWwDEN0A1rPyZHcnQBOaRjD49
Ltbn+hv+7keGDAaBPb32BElGXRaeYobw6JFUo8ylOhhf3tjAL+FIIRmSYk1RAWzvYS8nVGYjSimq
QfNOE7QGYQJY8Ot8/LnOtzl2IZ6llCtuW83iDKI1umzZlSQJY0vyc7GiNXLp1IVbo0C0vvaGGluS
jhkJMebIhAJM+zD0BEM15TM6jNelrW4wAnEiQ/ZNiizqMn2VMVimtkO8QzGB/ka3ta/JbNevncAl
pYCicVLKNYDwG3Ldbq9QyzzpayJJecpsz0hNjBobgu0I+wwg4tkB9MRqXbx4Xw5wwjqt6jOvT8Tj
cxAV4SCd8q6d2WZ0QH+d2aWckT4pMI+cttmpdZcbnD6gQ/8FqrsxsY7qW+OTjTWEGfA163S2MW6D
6UqdhJ1MIPFKD8be5eSfW/VB/q9wZH9TK2CmvSm6CY1QtGl8nR5+30pIyzzb/QsojTId6IpMHfJG
hvUKjbbKJO0iu/OZynJZX4aJCyX3LhlDrtVKSBCwGDaAd71AgmxDqbG8owT3bqqwtFodzeqjWamp
3DMyVYVKDR9NJNCfsF8Bdc31zA+5Ee3N5w2RkiV25EO0UsF1RV6nDGhKGz+EWnSJa1+ne+5gSvG2
Hc/VXXFCDSpNfqmPJzkzNamJ92YM7MJwehAlj0c4Slm9aasEbHPTyrlF9Zz5gk/QtEWuKVgVxRj7
e9NaV6sJpwOdY/rIkK2krSh/gcXIU53JZITh+qMo/d8Fmrro2W7CVtY7CuMFhbKM5vGvs7Kn038U
p1PPcskhCu0ozwIHRp/lDHrX6+kiV9G58hsCJUfFU0H+ye2KGu1dcAFDobxKjllyVwhoqN2pi3Um
3pwT9AN98ug5P6rXiYZgwJPhl4Wt6shnTsKejNun7Zj7vFj2BEhGCXMdSI8OTYEzg4MBic+NvV+H
Uzook3QhklbjnhjHhVESqBjvhfGr/9u6v1AUoW5yHjELQ70HFEDxDKdYcUTO8QscxMOI3FL3o81C
wudO5Z2epppg5JBR0OgQoQKoAPqioeZyjdYmjQRXGDyUDK2/+GSsYUwUxkbKvMw4s9kZmrhqeyx4
hGP1jglr39bb+9+j9IHTiAeYgOxnWmi21RvtAMUCsuAyoWXnVrLl0tvIjCPR76nmkbvRyQ8ERMYE
QpVCYvz1oVbxrfvshhEp+ArRGALYBQS1UA7LSWqLtns1V3bBKe9JFBvkaQDKF9GPeCZQpeNTpNF4
O81dEWNLMcVNx0MfGuNEigvNzjTWf6yT0HOKZPqnwr87XqCJp2T/SoOGjdDkITra20XIpqKpTM8e
gynqbTY6i4eyMozhk/G6nBBTGyoOvSHU5ux2iMaNNw4nr+YFwYB7ASdGaPFJq7sFxLGsNhGv8UOh
BlhQeuZdWsTa95bzmCQi3xXm9iyaQs6RgA1vXORAjo1OzYG8cr49q66sao38Is5dKP0HFdlx4iZj
hqjpkkpFrX0v2BoTy4Zd4WuNO1TabFF/xdAgCmVYb4VDbyBGm2poSTz38/deaz9Ia5cPObLvw/Kp
JSUjBnCY4WWbauE4KE22PkXrAY8WGbZ5u0cuQ6Fog7EC6PaOyR4PTxTp3UpEGTNPWjDi5Rz/rTKm
Ujdq03qY6pKi758V89B9Dsd0GEQuypQWSOLTfeBufeHR68EbGISewtRagrW5X2mGhRfhNJV8AcrR
nYg/xlCiwmw98mbdd0HsE88FhZfGootP4DWGaZ1cB2c6FvaRYWWFu0SiwuWqG4bY800rL9uBMQyw
LV/hTgS6cO7E9E1t9EVK+illTmMRrcbG6tyx8ELcXRESBye60hMvikRLzGHIgji4ClOAutBiQ+wl
gN+V/SuR843CCJdwZQzRC7RR2I/Ilw3WRdYBTQSsQ+a9Np4zM37STB/aEsNBU3yP+i92dn7VY37V
ggKMuN/+/ewxt1Zn9JcFfZYn7SfMPH0S1Okl36c0ykB5HsUTSkd7t88SQJT/SDg8w7pGK2pDHyje
zClY7xc37JaaqbQDcgSgPYefx87yI8j4w7ocGRQx8YIthj7c91TZuBoytBaAxTnjSOq6ffbIvTre
ts0BuJZBQ7DXFD8c0G3/92jqXr5nFuDonp1jap/Dryc/662eAw4ktFvxmf0dwSymR6yTasbMROBZ
+/m3hh1IMctPIJGqKSnUwRkFzKc9n4EUsyTTKq0GTIacPhqi07gKafntruVspsCet1fzCudvGJuB
hPI33LzkOJUaf9s9LfB051b8FoX6HDey6H8eoV18iJETSZdwyfGqCvN6chxs+BL+tBwl9vNcXywZ
5l5JYJsIOV2X1LOJEohAnGwIzsOR7uzlmkerdJ3DJHq3xGidoTZxp0XQgIYQQt3G9fMgxTd3C3v0
QWOPPe65i5jsVAAGIZ759gYEyimeIInjFtvSOo/WhUNvjO6qNdCaLk31tSHmLriXUCROfUvMuhzw
qcle/9VTaYX0yW1DuML9dAm0J+oPS2vci0VeqvQUjRV4cOob+s32mc3fmPGdGZnEWA6wjAdNLyP/
gJGsJjlX+uGyq26+vGYMbZFJEG2kv4wfoLR3wXnLHjsyq+nbtcXkHJmsYoEEJnjh0W6AUOlZXmTD
yZIHtT6JdPs8G4vvdR6jSLQPrnYkbmTy5pwxqJacgvnHs8hRan9cSU9YuYN0z0cn5g/ynqzMVK4D
9RqfXz2ipEk+6Ik19DJivbMgk+3mH9VyV4FE2ibzCnkCvMy9Z0QahOLf6BalXSeTASA37ZagxZmt
DBMSTiYWJ7S617pESgy/LyJnGYgZOWzfNT/cO7klb28pq/qBNJvQdxGXwRGBhgGcdsTEcU/b/l2E
PBJPXTiwK0chBiCtICAB3+ipO+s8HInWlJDTG7DtdsSjnQcWFYh9rrGKODBkovm8zM4YoXTZsRw5
rRjJkX5oJmylCciOW3JHjf6MqnaKD2RTsmNJFZek/uaLgaY/ZpD4ZWiRTb3jvCEps61v0X1Tpejq
55kXSEtcivf1I4z5YA1FSlcf6/JjpTFNGW+duGGlbpvu12OWwZXHRezZAn3tGMiZP+9c9ByQThJm
02cIlwi2MeRkqvYJBBnywRwXWd1l4k2jINPQCTY89BG9foOXys5aCFN1+aci21nRk9Xyaaj46M4y
Ak+VjmHahs20QHnO1LLs1PGMSxHwNQ3kDMHbztHXT+9/ffD1sw1gAjcwShQ+v+gsusiDMzXVR8yT
KNT8/PdUa8/mjYqlCRYuuIhqdxRXfumU0FezqWcfHubFwB7SWrJ1hveljW5YmnJTBoZuiAkQaZE2
6C6mZ7uiUi8o8cy4xy5FukXy6JlvDAgQneCR9czEiTcw9ZNTvi1zqJ8IPW7Lc91mIMAVnD2q4kH2
ra30ftxsUt9RaxIwKiAS3yjpdvWvN9Nc5i3Ge967jxfvOjzlK5SfZSaKnymlOPi3xh8MsYDUbG9e
rYVXLmALWRDVSAomZlFnKJYXtgcbtmhOYXtuVdSyco9J+f1bSQTEI1O97kGSqI1j7LX/3efp1Q9j
3raad+FhmBB8geWzo2h3pECf8y82TykIzPko2VAN72JP0xyhGf+RaXasj1MvsyBOl2o7EdXRlVUJ
9SA0beoShEdNh2B0afQQ9Lwl5ZVbe0KoaaAvsRJZGn8Nqyg0//9HZlYgmKMwp971IJY4QywnTdYs
wWLEykc2OnQYNGZhsbScE+i+Q+a1Ao6k/e4tCldymYFavAAkA++8qW7+pYvP4gUmJo76f4MNgmg/
6UfRhj0SsxHWSksGi3kuKQb8WUQZbBF4+RMFsDbdUYprpMyV5lwqlV1o/q+c9PHuNgV/nVVe4H8M
KPEG6ZsOiMi2D+v/kBzcNu6ek5VeN92tNWy2cX9ukCd710E6CqLYw/AoFvTMVtwy3NY5w3DEoDuB
tlGbavGqKpTx94S0w/aQJNxgwfCgp1VUisXEWG0lNTsnJlZ286EaDZInGHtq+6qmEowJ6yckmGvY
2x8i0zQ58kEhUs8/VIk7PCNuytmshOJayp+PiR3ioRQVJBJ5sX9jINIfG3/4bXB1BBJDIeTwCyCO
cZQUSAg1LTba0Epu6asgt8+hQ4A8KIMYQJyOuPawPhjQugyBDZDBPH75TanTiCN93TFL4UmR9hTr
63JwCi8zjMM8DxnFbS2ZroISOKzpEItirUKb6rz1Rqng7uiokNs9DeDUZUkeB0XbDpPLrLtGXWM0
Y+15x0azkfj1uV1EA5m8X26oM5d7bPrMkF915c/6ktTiIPH2H5SOt/OKh0R8H+OZh7CaGse53keH
hLMVScHvbMAQ57j8odGC9fRWsTepjC4LsAqzdLRC2HODG8py7G5BZH5TCUeQQ+UA5FKLIFBVhM51
E8jaBOFy3E5+XEGP7V+XJS7Yr2wd3rgrqkssK3UB22yfGgERmBkvCr6wWaItZLAKo+GodaqgvwCX
fF3YDEWI+MdIFaCS/lD+jeK/e5YBCk0uSK99un9L5abqcgehEM8AEbtJWssLyhi7sEY3ccaGK+3S
fJAke2UQYhzysPz1qzPpo2tFSL3cRu0O73j0FAHnAq2dEdqm0mvwvXXfK1RMMCYPPlIBriPqwzKi
vJPbFikE8G+ed1PRBfiSjrzyr+4EIy05oQBqZOUQuwX7uBWbh9qnhTZ7FwbsUEbkUxuL3q7OCLQM
rZoVeFMy7vq5X72RdsZXRW5ZFbCspQkWgOCFjSPHAo7QhdPNFRi41QA7JSIeCIUnivcaS2p1Afkd
wjW50fLUgJZC2cTbZpK67UfOlloy3qMNlbav6RRRAZ1k89/aIRtpd9BJn/tbYSSilDKVpWBGk5OV
OwcGgNEbUTvqtSgTirCRj/w7gxZxTyOFxw+qu+gmGFUq3AWnwAJO0iciWFkiVOS6q6is7jyP/HDf
tDvy83DlzsYdqBGumWdgMtWYCQJNXdx6dl1TRD11OnBI8rU1uaITzAUW4F+TTWDK+0cTfutkHGes
fFto6ZSzIoYOTCSrsTJOrD4Hgq1RoVpVf03NQNwiKlQC27s0mypqkJXyw/w+68vjvJDegfNJK2Ax
trC0XxgNhhe2thDrnhcl7zRdB6Vy0qcssNw7XM1VLRTq0VXvcviwDeofVYdERWc6OnbL4BWEQrFF
aTDRuNRwE1m9bCr1ztl4D4ru4rVB859/yGxZQoS7NhDq+QX+7xGkKpKW/LRdf54LpPodsde8L4oM
szrVX0QGEJ0MbRpn/XxXda7E0bRHxeqRqAlmtsQzt4mixpfHa/iBliawhSHe4nahjiZLwuBvO+IR
gCQAPzU8QfiHbhAFEwk2PUpyhusBEaW/B23qNO3tv1hR0WC4Xgo4cEtfFB2wDQI0Q7IixWs8Q8Cf
WziWPwD43WSwHpQuxdbmZ9zY430xtJEJLWn367ASwJ/wOb0Xrrmg3ILsQcm6VB9BMUR/InrIYrWY
rV4fUrN9wcaTkatUQVSx+cUovLuQjIbmTzLSzHI6q0eyz/3vUtXTqN2UQpEzThtTlkgmcbMuw+UO
bl2WPQ15EwX1B+c2ENwqQvZd2d2ysTdRaEZmMgI3bpYDMVSFF013xZBAdZJHQCmlMYPeac0Y9mav
6By9ZrG71FGTNJqh3eMEKvm6MlqR+dfzYtmTZxPneXWFdxRwQvn8EhJeaKr2ZmbQx4Gbkz3LCnoU
EYERQwXdX/B1ecy3wc05XRFLY1QZYG10qyuq7rEwFsg5t7DUQjWqRENQZWfXs8q5AVtTEIUz7Rb5
uGYBRsrqSy+Sehbmde6/MCNWd+cayHr/v/JnAYE5eggP8EfWEvBY5lTcmRbtC7rkapNQZzbvuTbY
bdP3aVYLL8di1f4imSWAqWOgq6wezkBPD1CFmQJyr9Sbx691+CaopGldOHn8c64pz9rq+qxvZULS
G9JuwE2+Zxrh6BXgVjreQIg33yiE9CilKdXKbQ6v1hlqCNg5EnlPBY3Hy+KSt7N8TzNMf1fA3KZx
rwIBc4wSx+tGy+iFTg9tw+8iN1l7qvv4JgredltljmnNIOTRzvYp+hr3skyihUaG86lwPrdLp1fn
8fKZ9HJ5GgxmI8XVVc6PgIbsxno5YspAJFoPpJVe4J/JBEhfVJULhly5KGUAa23ZqgRNTE0gIDEl
nrsOghwBfc2WFHGSXQ+zZxlTzbjnWTPsaUa9NJgYkBFfNlKOUUWLYqxCP1I25sXjk2n+fMiqEzeh
rrmYEnJO24Vh2Ck6hVwaVXtKIYHIV5Qibtp5mBMnl5u3+F2hXPlgAOyx+BjaqLHGIPnN82cC0aAJ
C1Gpu+C+N48MN6FTJjcUkcIddGMRi3Ragxf5n4vi7HpRbKgQJxNUrxn9LBLrbOp0d9la29389bkG
WKuSX4a/HWaEJ/wpbpzNKThegkgkJE57Bh9HlDd9eau3b/0b8UaEEr7llhLESqdx8qDl3jjPqR1T
xSSebph10pNKSrFpCVPPCW82tCfAxsm0+ONEMIDL1TlFyG9oXChwgoJK2nbYAGnB5d5I/KOuon7Q
/FHwBY1mUZu2Aamzy0NYFqK2D5VcKOokvhk04aRJBTtU1WjG9IVJ0OLq6t0IdtAizdDPmdSW7/De
81ngV7tri7gcM+K20iVdhlGdV317NLJjtEh8Wdc9LY3GVGa4oir5zJi6S1mubMxUFIDIaDtr71BI
h8eOFezIRlIYMyXDe5dyrP+Wt711r6ZZR/qSFVtzfHPaZJQcXZCKuNu3NNeVrWOM8Q3hnhTc33wv
Ugz7niXiCyaJEpqNCcTrJXtTKFAWIuEeUuosn3H0fT1T84cHGbDlhO3Mu1dUEJjP6ZACqO41Fuuw
kPzp3pqtlybfkXvviP1xb3glxD7IOPxUI7uuVED/bwLPxBOgXCzwSTqGu8hfvcJHb5WHywDxvygL
VvopULj8FZkAKaUIWySAAXgnfoi89ETjedwBqB8slW8WdH8ZXCnzy1O6x2b/bBU+wk/HyuIrBJ96
g/EmZKtyhWohBdOYLWAdt1uj6i/WP9UgEUbKBDB1+iCMEs9Ud/BJ3GM6jVH55IVB4R1OkoFmOdZx
JcU3Gpu1m8Ej4ApnrGrkt13WJMlnUctTCA4cxNBYRIDWHBqTdDRw1GikUu9krURF3B+7aXEo0YoT
XcA69j4j6bHLUajdT4+/KrXwo+UN3jfGW1rPkSE2wyhpoCM7S8eG4lYA545kF3kk/2KNLYuBp8fE
NT0M+YQI/OH9GMfz8x4ZF5cdv3DaoqcVRkiVGXxFXVtw0yhjHMAuI48nRtY2LusaaXIlEBdqTNbJ
Alfp/AWMnylqLP25pjZp5Xgsf6VZoIXIwj39mJgSVOEvkapyWqtLYr1E42S4Ne2Qtwm0s3R5N7QY
l/YKfSPLPkFRsm0pdgWfdx+8eE91oZdehjDpkCCLqBMEiys7WJGEvTzKlP7Ph/J1Q04ImaYwYtqR
JnaM+8x82D58l1AjzJG7LA4owNYpbVu2I4KIpsSzWXg2Qp/eU7vkJ/U0xGE2+ZMX9rdP7WZWh1Lf
c8ohCEuqJpflKJ6B4U3REZo5PCBYh9fR1QdrPqHd70GC6sy8in1q9KHv7crTFT7rEDo2zZBFgxDh
5OjBZbGaypZ2azGoNiiX6NYNljCVRbYvrKDlBMqXse8AbgwJSKpmeP4bHMu/vA7Pd2pgTeVtWL4Q
GqCED/lZnT1NB00En5i2QO22vG8FZneyFCk9rZTdEWvfz1VRnoqFW+EgceUI2/uDDWguC7fJkG9y
JDLuGeLGQBYkJVkAHEQHbPpXAdhrHSLVXkJUv9uvo9lUwEkpa9HY+CHoHC98f3HSY+yGHPHLoNTR
QiHZiwxvoDO3PWRzzJ17kfWwYhwJrqKmbBtHvd6A6tQxWp+5JLxL2pr3V+XZ5AmdXyDiR5Iq0iit
VwsDEjJiLppxE4obv+szEV/BtHO5wEUKW+2tdBu/qTVkyvX8znF58NS/3PZYtwUcXeQM0yD384ds
S0bPo8jyMl2VGwASmIAEoOurjsG2jo8CSFtRUQpHn787pAm2oXKR5rFAjXD5k2iOEx8DTCpb/5zs
4rVNSxpAZqzKaQAcD0l3hiKSdC9r7fzfD5g+yRNZJMIOCGklFZq15rX6s6+0Gf9n9N27GlN8b2O9
cUyn7Rt1LWKgXs/Rm3YFKGhGdzv7qNbWom7TNtg7thX5dT2nnswERy3aip8C/Uc3EnYzsIkcPnkt
cg6Krj7R35Pug6bx3VR79gszyDONVTfTgrG7wsAGOshC02+iGYoXAypPPUMEH1n3y6r75avEcce0
zgTQiGvINoFvoJL5Sh6VT2czB6jkDDChhUl7VGNWNfQKugEkN2PsPtN8IMcwx7etA+QPoHrgK69T
wl0P64yxlrcZSX59ZyiRBurKZMBUU3DTRhmTHgAvui77x2x47kryxpCqpXcTmmtQiKUCxeA2ETKq
uQyH6qxyEr4PXrR4GUb//Dni40cf3zTamqAh604aJm54WPDERyc/nOXWANCfQBRM+eXaDQej4Y+i
E99xfuyH6Q/m/lkuZDnTrYcsKyfuKRux003RHt8VoHyD9wHKUpHE+enK9zd2Ko0Lu6u/DzPoVJln
IH2jLmTDjldRDg/FAPmZBP2qgzMGjRX2OkqVYTS2ARWfAik2Dk2s1axlLhjVxqWuvgr/4plJoPnz
Hss7qWFVcyMjnC5inE7aEy+tE/dq6ciXe/BhaOX50ZSXnq2LGvXQCdJhsBLuf2TEm8ORkRa0Y7fi
LGrXWYFUdcFsQEPhZYp/3A9Wq73TMPY64bLpdBiUnRpzFiG5aNGBsi3ra0CiksTUiA2LA1P2E2VB
YpcKIKK9oLEqYINf3EfKki3RRIifOhOog2poAPvMOmNBW48lhOByFkpvrfB9ccE6KMSg2DQFP+Bm
7NaYpFM6aivFVaGljLz2nFnakuYpn3Vqg+AwGc5pQLWK/y/doLEkXemzogqyKZiPnnyH8qWHopvv
Vu9j16N9xMBw09aABs70fX47t877wvqKTJDqHMLqWLzkcWt7KNsmk/65RoyyGX39y6yR3zdcpjNQ
vPmk4IMSAdPR1PYqU7UZ1zfE99aZLq8+UgERcDSCWR+uXlR7I8/jFZLm9OiWyxIBJXQCK0WROOIo
ge31LXklTYQO54lJMEtTeO5KZsubUQSVEhksk03AHWdp6z/9Oz6Dj2bLPNd1bBW0hIxlxcUK+PGM
b/gyVXrMFDvcvCgQ/RwFTjvmQo/UaZ06reD1/mqVVLQwitKwUt6re7du6GivVYxd5yNzWhA5gdJV
Fz1uHe8wrkt+gvPay1VCWXPipwbm4pmRBf5ukLgZH4NcoxVxyff+t+Tf3206nDidnEiMCZrAaZeN
V6SnU/y5K3FODuZkPGi3cRvR3Hv3ZDBnRv1CwCKwqGbjLEKM/zlW8QZgy6uoDLWhkCIlYIdeUriP
mK2l0vqF9VCcUkBiA6xz5R/QZ7JyA3H44diwEEh5FPnYsfvqWPgexo0OxbX5jgOoktBs5tQHpy2z
vEGwZIxe2PJ0HfCjGgMpnlzaQDcKORKGbQAE1NEypGlpdgghaddH9WKVT4q8t5G50urQOOwYcCQL
BpvHnknZcUSTf816XUUZT8yOQR9197krYD0mt5D3/Vu8lf8DuIf16SjsRhANzOOifHZZoT2j/aTy
HgTSof97gZCLjE6F7dmfxxqNa9tP6EvRtwypENxy/36z6eHqPVf4zI11q/+4hfwKvs7o4gpu/YwI
2z0nnJUCLlUobZhN0d4tXRrvFtl8doP+RatGA+e99um/ZA+DvK0ACVJ8/9YyZbKrqIS1rPVaYVYp
V6ZHEqXm3RVkf5PX0XnpLnxBzdPkwVpnzqdBf4tY5Bg0BXwzGweI+DaQkzCT93snk9FVnzQGo5nv
rieLEPO7el+v0vVsvVOD6pjK8NqfCVLpPZwo/gb+sHdOtpuWzH/27XuOBd69ZRAL0LT1soAUVBPp
k/ON8P7hC/3cX5Un1OvTaOVllbsbiyuSe8jM9BgBysp3b5NZRLMTCLXlEF+RglmTmQdclLR9fHX1
0mY/cw9u0FMl0M8eNfYzK3C4t0+1/UBSj/zPbNE1L0DXvR3zHCvZhKDLpxI26Rn7Jhmj9hzp6bIQ
9J3hobUfGUDkLchx3F+Rr78rjEfrM55LASJANXvoMweyN56wwWUxnpVb8YxrxwHN6T+oyvdKjOHn
T+fijAPcGY63l0GHR1I/EgIIhqVX46V+gThvlRaVAEvqbKLyk+nNItSXDiCuhguw+DfK0P6OUc3l
V/hVv5RJj2KI8EIunNmK58/Vpeq8NDSoDM9cVuYJHRA+rloS+dGEfKuADr8JG7ohzp/sxToc/jV5
8ETQwceYTjVan71+As/71zVQwElZ4r7P5AEdVjH94HYiPvy9U0dRVLa7tvkk5GYc3o+h3N3fDthx
CwnBgF7zinH0Q4jGZ65WkdNE6nblh3ukhzlwpSKWjTbU33OUuRX9lvo0bMSljqOtQr9FcUEj/h/N
qZIVbOkuB4RIHKWp9yACysfWZEs7jDKnB9RIPV6WHm9lPIbCL05vduG2vg6obzIE6fIDhs3Zu1Gi
nn/4aL3hNA8n6l16Vpui7bCkvYOU7oANgxHx+14XpWnwGx+vAo7nsIeQApY15Y9ltSVmPUvD9bY0
WOkoKSMR9aLjeG4riSFhWw5kkScAilTzaKNvkVXNA7MKAaoMXbuwVnHaLr45NgfgLjDJV+RAx7Sf
akwRp8rcD3t8Oe+hmxTsBVlrt+zNHlfdsIRx2aG6wr7Ilv/QoWevxHCqtlxqkd9jLQIZdt/hqUjW
rTWQiOvYlpHir6zRyoXVIA8EqInIuAm0ZjsuujJPJ1q5JvHGJkONHuLxNzjwOvB5x7m0WisoetgE
gurO+EyOEBFGzB26aTIBymPcf9//79kXo5J3CAhSzA2Dk8ih47XIY3k0b+y4Rznw4Hb2jO8XtO7b
qI6e94bmgCUp/H8NbvvDR93Zigw7t4MrIsb/dgJFcESzZecl2jBcT7VqSvhwJJeyRgOle94NcLQN
5/A4srdMEOskRpCQvLfOTrRiXaBoUw6ztai326zE4WCDnIeFxvho3QSdymwxf/RZRx5I1f0wtNli
j8mVYRcg6Ir7Qprx7chiWJGbtiI5M4H5zXlxXt+JG4Rhzqg9IaTGLFlVjEKqEkWvQ8VG8B0h2Z5V
CGj0+7QHpWmCuA5Bd/jHJ5NEQdA/cNOyGPVZFuQmJPBa76TTrBUfizzMIXquAhsu++Y29VZAz5qy
BJfIpD8HpFfgqFW02giD39IuHJI73ZQxKluCPLL+C5GEi3Qt0xueEWyuEprU9TU2/2/WmrOVenpm
396de9IrkjUoq1aJtXPToz/KwyxLfAw6jA/MxDR90GpfdyM+7buU0dWufAvh/we+I2JwVf4uab3S
dcd5CXO/kY71zSIrBZfYQDS8MKjvMCuvJeQGOTd5RcYoPZ/jPLIXZleAMVyaBkeZP4T8HoB3a2i2
rD7Kb9raZMBA6fJIH9Hn/1/4JiDbeXuhGa6r1BC4Heqytp36U95yIQNpQMAvdAOXf+FAgColtsRo
XoV7cTsfPiVxGg5Qpqqwpsfifq0rjeD8wqHEuSjbH6d9uRXIA1AYPH02J5hukFJypa+igf9ejzWn
kDfE50v2tkxDC/Ap2ZJ4a0689j2bJwTS/KLf2ZrpfxioxxHvBAeePmNMPBoMJdPNLBVG/X2OowuQ
kmdFnKYMXLuq3+l7ZRrGo149DJmJcNE2O2U8sVYyUWx3wD1V4cTlYOJy5CcjOtS6/KekKDEJ9XJL
qPUI1n5nQ2NK9vba+WYE6Z0g/mLeNqNXNfgO6ZGreI0F/UXiOmVLmnz56Nx+G5pPDA/A20PjdCxQ
tIVfIlUp7sTqoeeIxlUofz2Z+gSoVFeAcB+ev5gvh6R1f1P+/aUFrnq498dMtAdMk/KSyWj9QDzM
6Q1YdKCf9IL2JMk+w3hoGb3jotSZseLOjUdSNUs1Ozh5e/lpMEtmhIfBaTClblEVeLf4AYc5slF3
N5LVB9wupi+HuDEOcKFvJt22KEVsqiwOaVVlUOEjPkvQcYVsBhYJl6BqySsh3hvIt/52wYc+1ekN
qqfwQ8iVb3cFufOyuVcm5GT4UqgOMcBHkG/sCu74H2baY6Nx3KeXufdFq6kRZ2V7J0gYGxo1jNtY
LXoBuaOTnynH6G2qxAvIwhdrj2cFR+w8Wblai6QdW+xgUsAENZ8YPdMWpKcPNFOgLhohGHqBZAr4
ddEyT8hu2anxG3iefZqdNcmLR4pr3YAm881YFEFxp2xASVGEHCMBRR5E9cjE2AGlit/LYspEfuI1
v61x/ml5MsvNmiXmTJK9+q78gAMrfInoDUjspjruCr4oPChbSb8ghy4ItVeMhhAqoEyCUlTtS6ee
q2vTj1AiDt2VF9HErUW+ZoGJFaE34rGU6YJE63ORODzbhSaES5adnQqLFtIiWEkVb9rHMlKG2Yt5
j9gX591w+N2OHWkPiHjopg1Uh0JG4ZyZfQEBHAOJDMkhblISiaBUgpyl5eqz2dXzfw6xaz4lMCl7
+gSbIVTp158LkoidzlLegwrdyKBrmaaJn5J49LGjie+F8uQAhKQpOeE4QBFXR/g1S8xgxn+Ei8lF
cjoM6SA3uiiDLG4z/s+ieOhiwNaDbQYu8C8LTxFevJkN5AzXJY4bOiKjlHAXVG+JrvZoKrF7Q1LJ
DdDzumGE+py6chp8Rx1rsOZ/ViO6AxPv8JmBtVuLtFBwzaZOL3xFN2l2I9vDkQ21Svf6TxJowl0s
dg0hQ5cwFkUB7hlTdYxe8osCURGtWt8IzDjLDNuwjK/bFjMQ+cKaVHAnEQHTUlpNbq40WbxsV4u2
Zl8wKgSjnTa38/j2JGqt4+ylenD/gLQYuP7j8ERMtV9477WPBiT9io1VYqvmnZxK0LjLpInfKlxE
iimo3lQam9VMURpcVmrssJw5knjjJZGrTThBsPz4Wjbfq74eWxvN0qcWwR5KuqbBTIN1Yb5DJb+O
+nGltdWETfMpAB5N46ZVRFPITVRRjmWYu6bX77a4lKmKmj910RhNPOUtCuBMqaCvneNpLjUCgsvY
oXqojsaYYZTtgjY0TLYu99bYNMq18+dyIMysBWZGHq6F/gn00JmqqltlOhL5KAtcVBF0MiYLkEi0
GFj7cjtsjTFenV6cnPsILR/+V+SnWf/OwRzKwxvz7lc0MvDtBIsmW/Wb+u1snCo9H/1CbstsyME3
iwOeUxU+jgCpnmKpG5EhWgzBdqnEdwRIAJyRDDShblaAHj32RhEltbhGIICdFz0zb7mF+PfdpSUI
xgu0GcZxYxbyVKuuVNNKBLSE2l9Dp5xivWDX26ARtNpB49haaH0nKmE+UxZUdxDEUv+qNXFAK31L
rKaKJhuQzT1hLyAiA21Kf8ldm87DJGT0ZOnSvugeE+t5qHVidhQpq95q6OvZdbh3P52yl2hPwjvH
O4omkmjmC+iaOcRlLIDK17ln/ffXKPH8n0KdqdHYhHoerzmQiPnqDqHF1oouLiKdAtVvGonyJ0nj
5ifyQ+I1Se+tMRTAte6msaPNWgfT2mdDFygcViD3hY1UYkRJbBA86d7JKnC82wuj03w/sYRQucLf
ieR7SSWL3MpgRQ/0ZGYqa9aaKSNWAdDHzA2THpexnDGGR2VUIZEunmmc9nyWUaqfwkg7RB213Hp6
W+pdMcHmpE18WFQqm3yz8iU8bxJBvQyVmUxpBgKfPhsmmUrgHAvk36896j/5vV9BCfjqKXku65J5
Zi9iGmgSPyTPZtVNp2bHuoRQ31AiWCZCaz5sZiVLywdPMfnIGBXYclCOYBbXbvORiYguzXrHkkhN
3ygUNuolF3Jz7Cbr4bkagdxcBzayHz4xDe1tyv6fTHhqh48glmOXblmh+P84eqrmsoZZoEDySnjT
Lw2ZyzAoDG+GEGpToyjtwcKqh7gawPqiQSIshwgIeS6E5My/1hYOwCEgwQeQ/1yM7ZdiXfQHAd//
qJgjkIRJSDQTY+tcUVU9uZPRqxbnm3MsWLlr6K+UH4kzzW98g3w5my56a3vkOuVVIvBDapbj9UVi
gdjpAk3+GxCrcYsgtI1ngD2WpS8PifThkN4CSpPw4KVB0UJm9WO89AjJbNRtBgVmZDWkvUVQRw6H
i3q4vobceI3VNDuL/iPl2HQjMxfz6ZoO+7kgIOH03jCKyhoOHLCR0z6PURQ4i1f4kw+EXL0qvQKe
ycAuMIz/diPXChJDBcZPMGc37SrgxRZp0DK9BE39lRcGQcBpBNQB2SsB8FGxm1IN1UluwjQdeHw0
8GECUs1AcNJFf8Xn/MJ3CRKXCUSofp4/mMjb1IB9pfYyd86qDJjRopS8xe+Cgept+RXc6gqUF4fA
4t95MoFpiZp4l509B84dsQMmImEj9zBvUEnyPlkcDxqUGi3j+E2qg2UmtCvFBj0g9p8Z4TlcROU2
LTOgYL5/JnMw/F0Jh0sWoofTMrFg8hV+S1xkWETWhoeq//Z1fV2DxsoEv4NcB27ii36VpuUBVfIZ
gPltkd59/0kUhH09UZAQDxrDWJ9kWLx0ylRvv2ezOmoMNrLsHckD+I3Oof39aHjhyjzkMLiVDH1P
XLMvicZbBRw+0O8qWd56/2aQIjWeE67w3YFNbqZdynwvGH106EubBIpMn3K54VKU95UNe9vQGmJs
8NtvHuBVLPdNOthwpMSqi0SBnpVGTl3EeS7Jz7JAhmAx7VxUq2BJW4HHP6iiXlRvCs1TGJmM398U
HayA/TWAsebl6W5RlGW+jeP+nUyetdl9Etu4qq9IToKqe9zyl8nfr8PzkEfIge3fMs4uklUzIMvW
LBC25ADlcWn3esNfIDNMtlQ3kWPY1KMrCz9LrNIRNsBcEkFe2ftGAWr3BsjwmF+WH1iSNID926vz
5VgqHDhX11wuf3HUPwVXoPho6RJqorwmhCCX7rLEzGoEQjRUB3J06aO+2iRN5YvJvGcOCEm86jmp
hshwFBYgZGi3abmXUm/evAbbym0NZrY2Rcg9suxp5I5Gld6+oLHF++ALbxa6Ziy2GccNDYCwvrx8
yS9uffT76T8cadFzQZEJKm2L+VNT/tu9uhEeJUvOyK20Z0iAkJ/d+NlreMVNdpZjffqG6tL8m4HZ
s8bv7fPxM5geD+GlQZt4z3f4lEaDhREe7C0JY2NyS/IxwtWplF2h6tiA0+aWwChOsGRUMmREn9x3
OS7OKfPT2AfZwaKzE83+N3dovCsn/xaBKFlU1YijrJV9sa19FxTHgm0+d6P2pQ2KM6IugsNktsSA
uL3S4MEhkqOUptYol0O6T8x28SnzbABOWxRPTUNlnK9NrDIGtrm4OHK0q99zi6KI9A0WJGqtsH3n
e5OsTmsQ8Pcoxn2vMl3QTiQ8qNOVk3/EbY91F9rPhpeiE9HrB4cF+ySv9OgvwghWyI6mpiwqKPqo
56TuDNoAHBtJahJAJQt9fhUI/Ph4DWhnVShweyDJ04njWMUzJABRlLQzsJ85kZBqdGBN6lkQqCYc
OjtAYPepLXNUIZdXPabAmNR1W5r8Ii55bFpnoJmrJdRYklD7vZ6C6e97ow3OB5YVCgrlYzZUmquY
2OF+CtB9SwvSC9tzuSzZTlUgo3nxCtUYW52ngQId7EsmvSBKnr8PaaBA6r9qvOLrKySgOdJaq+pd
up/jmIazTKe9qY06n8OvUEIxG56+ikA74zO/yyLagOmWrmNFyvUJdBmpO6CPM5MkxOZ+WIkXphbp
xCRxl0Y3ydVJ2P2MIadVIbiaV5pH9OJIxzTo7E0MJLutsYdbO9fipBwjqIUE81LZTlaewHalQDkT
qdWk3/qUSNPwJI4hheDV/ZRDy+GIpyXbzuI5kcuYZDCzaHjQ9MjS7MoMAuT4JXaTBKfbdbVjMj9x
IxmWl+YWFzLhOaC7rb8RFYtGuSBrAJi5pgo0JbZtVFJ2UC0up58XiX3JCvnSidIrJ5wrCVV/JZKs
ELKSvDOLBq/laALdV5JJGkMUtW1SOigEapc+Y4gG+8bqUT7B1iVbOZLlrZ4erUtnWmxz/IjJYpHz
EOw9ku596nC4XiRhdKnbAJvFrSZx8u+LwQb1Z3hrtgX6VsUqTisZ1+N0zPJLa12CXmmG32ZeZuC/
op0Z9fS6dVt9cM7yq0h0EIqknEYz8gKMxNNxjGrmI6HrlKCCt1Pb94a0mKPNl0mjGzLABTxK+x4G
gss5hI1ilDqXKAnxt3IetpYNDo5OVeODsSaTScimo8l7lA02ThQa2cC68Vlbei5OUoWGqu356VIB
fXh/uqv02Dfr2Lr4Z0Dpkuzctqzda/KrMfNeBJaM/CVn1nWGpWEnNwzx+2M9gePvBH4BdSDc4xSH
qcuE0SUAo1bbHaWR+XSV/Zvx/F+SFHqm+nDLbtWmztwiSTD2+mZH93gktIGFy1nGHJXRdZibXTKA
ywWowzAvYyNYkqpDM7pLw3gnqXSGp6al12XAktq1ZML3OWJKwY9JkfbNXYrTXdBpxPSbcPqR8b7p
BCUWmb6G01xTzh3STKmeB6Auf+82KJ0/CmCm2a/BmQfNvH3qDIL65TuE6lZ12LRV44XwxqXa0Sli
PJWQnVo0KCR1CF7A2ZFayaHxFXQRJRCfuB1LJAh6uG46nQECeddQCL7ri/hpry7sEK76wXCLdZun
PxnUZWf1i5YaGgM07ou5KiZQ+dvQRkdgMkgkydvZmaiaKsdO8OhJJ6AheizwcdMefn53Y/tiDlmE
Fb3cRvrTzL3/F8bp4x9PhlF8RWcWl/h3KCs++HuaTfMJ4pjlogUJ6hUPjbRvla7v3oIRSm/Q72N3
XS/kTo7oSSZZdWVqcQx8uy3quqs4e0tFqjBD4xRSfkdib0dwreICMoK9kY7rfPRpdd+uj6810CUa
UL4yqZjTD0HiSkCH5cvl9VFKd+S3scuVm3ATRr1J9wXnfdB9LfbLcK9Uiuu9525iAT1drXCxOWEg
bqiAzf6YvixZRX/190ni09Hfxt4ioTQ4bUowFZHyZBJEqOl3z9D0v92vgl6oO7PCcq3q2lCAhPWu
UqbJEjINMUxwMVV3gDw/MCi/2cCOPwEcP6ylUx5+n9DGKvOTE3Cuv/ldFEU5m526rYOME5D2IlOw
/6SkZyOF+/Q+TejYVf0uHAWJBgU444CLqVUoH8+EUFA9hTrLIPsphEql2435PoTtCBNx13NZme4B
8gN0atAesMDVwkzuIPCfeR+yZaPxdjLPMkUrs/seYits8IiBvvy8vixe0Qb8ml4NTB/U+InXtYvb
izAxn1Bb+o6+6T5GZfiI3Jg1/cRWo7F1uAYH/Z39efdq7RKLqr50gPsMa1P6VEGLe7KLBIERX08H
iwh/jZD4FcdtqVadlAcJ5VKeE5mTZaBavrEu+ssnrTqFPhdk16KqqIitpaoe8gQTgCzFhzEuP8hD
dQd59mQQORotgFLX1KQJhuOKR/NYwn8411LtGns88Bm7wClMl7ARzGgxO1859h0G/WDdFVg/3984
1OrVaJ/62egAaBPnZAI1hSr5ngwsBo7KPiLAiubSUOoMhETDWlztTmQmrFe8hscvadQDORO3UBGS
8hcVigVVToqQahq7BsP8RAT8PzEjLUpc/HxAHpGXynLYc+oQ2nNLpWXNEGcWbtNFC4pqmDvx8h9j
/oDncczAOn66J6bh82Yz+PWLffNR+VjcVj3yosHLQ+SJOuyVx+kbggQyyWPuKePNJxmAj8Om8/y9
VTKmP2YfwKlOP+0NNUAXM27M2oN3zGmflSj/b747FFi2G6CoE0thyPphN/M7vv2VWpu/ECemriMI
CHs+UEN4hg59m/jJzIWI9t233Am4uvEMXV8ATtGZ5zgQCVv1WCNf4K8r7HSrP/XzOrYRnzGtcRR9
ERH1mWpnog8AORhBpWDIPGWAjLhBwju1LMgLqXpBXUjr+BY3vCbwN43kbqO7N+bkJ4mg5iadWATQ
STfSRILz4pfGT/3NFX+gp352B8GYH6oj59dY/xf3sEtpu8wtHvIIQB4GJBEDPvFxgyL9+m80kpB3
umrkXD0m3TpV8DE3q9R0LLoR9IZPqZwV+Y7IFohXu8dJRuSd5sCFnCtTBYE+H70RuuEFh9arOquR
n+uEMIfyLo+vdbuI0bijdksh+tJWm+Q6b4unHQhHOCUedCUhnta7KoNd/lusv98WqcsM5xsu2jKu
XLxmI9wWnW1jJgX7uMjcCGLPtoYHaYs9MXTHSyGDuwI1DrWiS/d8QTMAoUaLajb1CwH+EldVgD0r
d2RkfjEHI6N59AftDR4/Zudu8HvGVsIjEf94isvbXVtB/IYtZKnvkTUd8Hqup2KmxiVEMTy/2upO
YXxXFVRhaICtQziR/Ufwoe59pX8hQVoiftclYMOptoGvopnV07+mrjlbCHRhRPtZ84UQYcYw91h0
V/BJe/ugA0NsJLs54l9INLURAI3Lvhm67JMjZ/sfrNJBtqFlxZkdkdaDJEbHDAfvr6piTmJv0W7n
Nc3Y8t/3l3phxd0b+87mLdQiz/e4fU4gn37HySOgxhyklZiZy7RJAgM+W4UHA2jBXLiqGSoo0BXw
cpD/56WoqzW1S51EtXdnpbeOoqCD/GReib1xAve2W8LXloIH8oKCS+4q7x8FNTSqcdL87cirvemJ
5Nx/wzSwgEsA/KmZIj+6nXCYgXrw9gjpSCEfnUMJKiNOnvQPPKS+KJ8E2LbyjB5xzWSaYT+LwBIn
/Nvzanvxf7ioTgoT7vH8g5I6wXrp6mA3M8ezDJnnaIM16uVf7GhawtqY1ZNScCAaBLBxXLPff5xo
e2aXtkzrq8FPkW7N7q2hbjvvsP0jhTcPYwqFzb3jAOneGkdClKFmv3hj/dd8GOcKsun6y7JV1dJL
oFjGMuBoSpm+kYdfqblR7LxFLf+D/RyRUc8JGwlG1kqAW+4f3VfQiH6EIa3nDBQXi2VLEZVhBSJ6
adt+1jcxzvFF310iY6EbxS2PcXA3Y53VDj2PPGUXeqRBVYwNoilGOszK/KdKKgsTq7BJV1H8Z3ZR
io8R2muACiSXU+G/DZL/mTMbV3YQfx7l23nVlGZcKs30VnBAZdsO8hWgWWKx0k10J3+mrq9LU3Op
hs91ZG6epq1LyEg6SoDlJVAmsG/yeoNPc4C/c5LReS9mBuEyM7eXgI9VvKDWv4pD7dzpjI92vBQw
5UV1am5ZrxnJk5ttB8ocQ6yAw2sPrX1t+eC2t8Pa8I2mpHpYsImtWvTxe0ezi9xWVgp5pSpxhynH
I960FOx0B4viKWiom4etrWwqIU030rDUY/9WBkScFrdmhzvFxv1gCMaYrqWHcqR/afnUsyBN68ux
3kWV7Ifs3J+DqGXUoZ96QyKLm46JmrtEfj1FiE+/FgAwHyeJSSa86xY4IIvrTPyK/mzL5zcbSEYK
xjwDFpgfncACyD5LYxDpDoJ+J/RnZLGK3JAmq+xgOx7HIGPNyIAh7gtwG3Cq4bv/KyaRV1WbQE+i
5EQYwF1Qro+EUuHMLgJplkp4RY41y+6gGk9VcyVmiUV+V5SNp3Pc4x9RFC7ZQoCc2q1tKvp2RVyX
uECaHu7ONzPs2G9TmMlwJraxlw9tztWFYP+Jjfc8fsTsHKtIz/I1adrgaeZEvjxlNcLQEy73tiJ7
OoZ2+iQJOSbUsZHpLpPYhu/ETqDQZ0U6wp+lbmmpTUiFV3+SwAdxPQVD+qm4syekh8/iL3a78svq
48TYfFCNCRqlEIqkN2DTcEqat10NvXzgtMS+5resJYWPM1NhmJRmhkg7fM7cLIQUgXBqc52Fmwlh
CTAk2XjRUvIxmEvZzShdhdLdF9gfNetnLUD9nnU/D3wkQ9l6Ro1hQMdYosKGRxfVk8BLAC+z/VlD
wuJ/PYn1TZ4aGnoAY+ppplKsqIwOVx3aBFbu4y+a2GBIKdNmewhmlGw4gV9tw9IEEuz7xsM0Uu/1
GJePYMwCSplDmcAHcMY3DLmb5/rvPf0szWEtXlFIjPnA0Ibt7auMv20vfBtNy5yoTtRCgM8ehEkb
NW4nP3dfTi80LvLlHwZcaWU1avLCELY+LTeII+75i7RtgDcsSJojTncL/YQTFHciQKUmWi4YrpAa
z/5ArXvctR9TIvdDowCtMz9mZBrsn0oiuBWHyA52pijlMUVhQr/Duq1hoQDxCYj0tZR18epWdwUl
rSXrn+xJovsEjzerqYXrbJQ7NyYi3THP1/nS1tccs6LrhAbPUsxZ3jC5H596Lg/9ojp3bD0eSLDC
DIomAe9zhgz1wPFZgoSlxrA20dKaU5HoslsfThbxlOqMbwRYehtDlhby2icy12yp7pQuG4BKcJSJ
7/G3b0ZRmUVOjyr9ED72qpEie1l6tfLn6JcBzqMjx1afydF1u59AtnOx+oI7Oq78rN0o0miqb++O
Q3HbW84oNb8HsAekg6J9anxarePVADA4P5gyIhG+ir+4AKlP7nEG3eRiJ2s9h5IWCsO1v28BGjK3
Cd/SkxlaDYSf9il4gH0bUAe4/uQnwtqrhSyynE6MzrnKHAtl2DphaKA7tWKbbRW/OaIo3yQtuT2a
dvFpXJD/YSswOBzyYkbsadehnWpPEFAoAD3cdNU/wCXzGKRJ1945C489jwdy9PaMQq9DfSaf3O+d
8FgNqxzUs6R6YxZ/Cl6RLZjR8eOXrzJpA3BFZwOV6A9zOKyLVJeqNZdIJyM8+lqcDK8ggTKeYOBJ
xABK/jfkvBT0kC9TTcdxyZ3RCTYwBWFg6XakYHq8ntne9CgVhC/4pWQmh9jqUJwCSKufw2y7i9Cx
MOqG0d5tI4hOtvWfMV9juQPyCOA6dP6kpQy3L0v4IgZILIwfPiywVz4j3ADs0BVlZu3OjHuSm7gI
sPHdqA8+GtVcr7ztBWyYlmkD4VMwnF01CmapCu5UkQXjBIi3jtdRsa9xSsGNtXuspYT5pKYWY80w
n/aKr/ocKL1YFHPyTP18nt92nN0hXqYWvgEg4ZOzwA7zxfrASciUarQmQ7CjKMYwIw5cimvpqNQ4
KasnQNDR0P78sHLHP3IG+FjRgDElL+5p8hv7/k1Rwm7k9r3Hn3o6Nny1lWiomoFNY02oUPFCf3dD
vpnX1Ti08tcRlk65/qxggUKUrOYAnW4hudWIqUbRPuSXpVjvBI5TZI68r+RS0tHBRhe97mrH7W4u
afRrK95VLq/9KUGKGkzuuv+W2l7x4R1wn1M8xaLx3QTIPHndC1d6Kb/45BiKevy4qapip+RTLv9r
lqVfzjyWu0/iheHhL3Ku5MJg0jNfkayrA/L8O779id1URo/JYB8wbMitW1expda1fwN48tQZO0w1
RvCKit1ix0wPsXgQpfMIxG0fsREnKgxgQDVjkYgpiYkYgyfn4j6HUjC1VYL1EzWW0P4UbAemkhyl
wRqi9Nf0Jp1E+1kME9vow+ovfLgBwXDgISJpD93ZWVYprlfdUVVEBgREJrhIIQCAYHh23IsE4VXS
7bjm1jAK1W504Vhj9vBWipM0//EBdbcmnYO4ZuRWuy3FyDQAOpRvGtd1DWyOZaMS7vj+/Kix+wss
phTn+5z/zzE1qHAJ9I01vNlYmHNrtGpPwcRYvzeYebBoqufpylM15mjF+BbEP7sYUmRjwiDzjA3e
CtzGrNaD8Xosbbs0mA32ZlXwFb/MznR30C6GQWG5cBy+KnST82KB95Z2Jji7eetnyvmTPU2b/hnL
z1re/+vxj5SjWnjrDrDv9Nl9GgL2HOCNohX60Z73B7nPVxRFEgQcy0RAs7izRK9Ti/UP3Yu7DVNj
DgLYwVzPA+miPE255meHR4RzcTEPEeDaFmTVfQVlTwdsEkrLH1JunhzJb33y9FLq2l80ViZ/4zNZ
FQYHIdeGqggFXdLH/zunDHbhun1NDiwqy1JQI98FQXwPIriY/0qjEsk3gslF0MbHmaKmVZOsTIBv
EOR9dv7jwycPUyk2tMFJhPRdwGcuu/Ve9a2JlqLqaE3RosM7VASpT/lfG25io4AOIu1aniej/Cgz
5qg85atq2cdhZAsEoVavq5pGgoKbcHWpndeRg5dRY155tGLKfPumCo/0z1Vf1NqTOpS+Voa94oDe
MRJUNTW1eRRE83Y9IXzufQkPwWu2Fv4pSIoRu/94s1ZDVBWn/9uGwMTdzZZSLMFJ7Ahks9wwauoH
ULIPe754yjiWvNOpOEtcxEm0h56owI1YI4KJzJX88EB4AOUSfSVM0UtOt11QHRw6bZdiSl0Efngq
0lH99ZNMoF+MsU68V1BC34i5SoUo9uGCaIsE5qmiDfxtg87BL6m0DfiWOsCe+LmfR934QDONSZE9
jdETxYn9X/gQUjdI6XE0K3wRuHrU/15rMUGQiEZKwUaVKOfl2FVqmVMsVfyufdRQ6YbONyWeK6gn
opjFjcQAZd+KsbJSaF2inkVpsofYbprVIvosbUiAoVBxJgsF477FICYe134khIFr3pSZBz9Jfa1f
oTXmDmhzkXcBIl++KwJQM/PUprs5W3VUh+F59WJWqNjmWNXsHWxr17zXBgFtBIzB/GhS0ybko0Fp
p9HxBE/U0r/oIlCrOM/aKJiI+AXer5QJ5Rxry0s0OKvVotHsF4afpb+Cix1szPKMPHW62qLgT3e/
5Mm5JUtUzWn5YCkNBj/8Jcw4coYySfCAqn8yy0Q2WItMYEZRFUMxuIy7VSu+iAM601jgp4dDcd5e
Ew7U1Q1LrcumoGvDNDUPcS4OqmKgfiXm1dTPW/bSueZ9I3IV4jVEBVh8dcabRi4j0TuWyj19xokl
xaKsHuMKf877QhxR7/4LqY51o+NYlf9sOCgpXegaLy4w8FdPJdImqj96cVuvm2mnyJqNuRTTAWpx
8RLabtjzk7ztihWJLruhip8397DxSUKccUZd4TXoctLCYJd5le7FNDLUY5cDj5OB9oTdewft01BI
1ZQJONEfHwBxskh7VLM4DxzqWlCo/4NLZLfv8s/guMPAr5HjNQwFr85QNeXr20YAj3fGuAHFa/zM
UMLd3c/zCJzeaQWsE1iOPJfovW+geY+42oEw5GviUqPFm0zSnckzkfnft0ChcpknihED3bC1yt10
17ctqOPKb/FeeqmG+Vsumtc2bE1XKiyy5Mc2/UauKcwnYg5+Xq0qp5yfFJmSL5EiXnj0i3I3WzbA
pwGD6V859GNjJ64I/SlKZSB0/h/fRE/goTNxb+53sHGYOhslWfYeQRtbkuzatFYcatBM0PAgAqxX
lLM3i2gv08nmVraPHgUNJj3KVjI2bV0HYAzeByq5GXpDavn3Y95wIUBtSiB6HL++SjPQuAMPSnRo
DufWzca2JXU3gRT8aci/waJGCd/n7+DCHoTJ4l1nx7KR20iTM1FXmg779dRDFmYJHB3dkI1KlNRd
2xPz1sN2+p1vLJwuFvXFrTjV1LysYMcqMgOYUmML7XIlc+xNa97LzesDhTNPQ08PYOR0KPvjrp4W
1wIUd9rjSESCnaMASe4+BebgK5/+yDGHweYSRFINDdDTv7NMplcVhSPlFnm0iUgSIAGISjuMIAl+
NYbQS0uthmC0mfW2bnwJp3+w5NqKCiyJWW8JjsVpA0unpXq5qZc4YlqolCsyJ93RlpGOeT2KNDEy
V5PlDbOBRtfK9pMZOqpXxVh+Zb8RIVfnghe0D7fKnlZ3YYIwJXBvcN8QTE5H+QDXT/EUvKJpCRqv
79vTF5KrOAZ0C72WoYZo3hI4Sg11xuIql00IeBTVRvF9T0m6Rf52Gi6vEakiMnuELLVbaFWhEoTK
A0CzJEyBMUVcXxcU8XlyBaSDYuEWXW98Gyu84CODB886qh5YvDrWIbMqY0W3BVQAoYjWjBUnnjmY
CRKd1m7ynu+hZeczC8mx/HtUI18xp2AbA7509WwPFkV7Q/cZKPrNF+9n8J+d86Vl7OKpeN8eLZMh
l1dRMdVogVpbe6LYOdn9/pc1lvOXOSLs4xdWIzpn70T7GCQor69U5ZkQL7GJNZyRVqq43SfJVsI+
BWSPbEiQgLboqIV0CoiAoFvKrUfvZEbee+s1nHT15grB2OA+4Yj+GJMbR1ztFl3V56ko/Em6UPXp
oRAFJNZ62ifPbabnSSInXdV332t36rIfaoMR1AmDsOR13oHt561kKHWqs3p+fXzjjDrUHJIXYQDL
OjCDwRhgOc9wbWNEfnXRuRHio2FpHVtMvGHwXeu5x65vYmoxvBU1V2wqkTJBEXlhSOJ2fImyWkRi
lRzpAWYB6UYbtwMcLOq6RNfNu5qvBKPOszitsyPU0ge2uEayB03a6vF/bwqdLfqbGAOJPPGUcu3G
hP/hZVcyLqBigavaZoGaet7Gmq0fIEWiu491mHIGUz6RKSNWQM5kD5uZrGZFUdH8izbtodz2UR/b
7CQ0+nSUW7Ukdf8tnsw33KSw/yOWLzwsMcfU001fPr2CfNNTI00NJmYxa4c+GZZXchjOjA4ymzPU
ofFmAteCe8dHjauM2HAT3al/yMMMOtFIWigyarv/u/n/Zsk0s4rOWwEp3HMpigRnFETo7y5WRqKz
Y0tJG25/RZceJ1pmZWUSFrm6YuvRj4qRnhrzlBU1Uq6FW36XSRjQZueptOTNDtZNWgqFa6g3LiMn
aXWQK5n8/rngZXtuL6QKPhSG1IU+siv7pwzCs8vhs8cTPD/Lmj6s/eGSdbcUKXXOKsUmFs37MZcs
+wxUWw3Ac7r1jupkvuoXRH8Hm5YWo6XV4zQmPqrp5SptE7h2jnkLQlJ4nPcvZbOZ1rbs4m3paGCS
F1wgApcrJVE+g9KWoxxC/rayXf0AKoqwvitFCRVzpitcoECHvSxYttMeKiywXGfYxPv/tQeq/ruo
PI1lcLa5/dzVhnsWN4LUzGTaYPXrHiTX6e3E03/w/lLT1TJMjScUm9yq/csNXmJXIWkvGG1DxdDg
DUXk1z7WJ0ZrddHfq9HZQ3o5PO9wjkIFRlQuMkiDuPtai2Btrj0M84cKuvecY9qAD5Q81MyWQ/o9
hVS7EBqDwf04P1sXOtZChdDvIbNKGlRCsdszD55ssfFqCAyrJxdAjBy/Ta1YgBACjQ6cYXV9e2Oh
lFo3/51PulhylKPX14HULxbgX0/EISsW/EsSdNtiss0sKD3wIttNzFWYiqTxxrAvbcskDCuGc3yQ
hl8yukug7yuMyvynGxq2xaV9iZEU3m5GxlFtvUZi1umriUWoUog5bPWwUwEb9gjQFAIRvbVqQQ7p
IhdEUCICNehkFBqEbBiJ1ySk/awAN5wl7tRL1QrfDx38ublOxTa2VnBH6ulHdfaJ2YqRzB7IWrMy
H+XMpis04Mt7nxXGnG+ynPhYHa0noNk1qYTNz3EePKlw+X1sSGZV7hxADMVJAgxNr4mBmPAOA7JT
pxfn4sh4Q8zhk5tX+ffMhw31Qdpfj27XZaBqFK+ZB6krpneMSynygEveTZEnneKV0PYV3dfzw3Mr
RkQvQQCKrM92eNsKVglyfzkuflrE1WR7oiUsbfoJF5SNh3XcD0OfjKtKEpIGEi8J3CQcZFu4Z3p+
NMzcdnuQOaMS9g+KLk2Q18iSCGrplXxbA4Q6lgndynkPBlZ7nm75Y15BqlBGSOhXEqrMOidO9DdS
NWP4q2BdgfOR1P2b0slq/R2O5hFuQqnagnbmlbToJmRWWRTAdcE0kL7s2wrnqtsMXtKGF1yNwQ7K
e6jqXUWg1uks7u/eUrDEi8vbS5xYhGKwNAjwnZGO3GTwD35N/CxIiM86i0zRsZn6Lat6aSThhfxd
QmV/lT4Va8DJjINTAMBJKNHdzmsCf5a3D2StXLEwZE/ZyEsfCbM6ptkzC8wu/vBVCGTxba4zn2zE
ndE/DfxYudBkba/7VsGW8qujMlj1lxc5L4XPE02/taArAchH7+EhY/oz1hwp+41Cm4FzDs9v86Du
EE+YZc6QG3iUjBCoZNWUWW1asi7v9wkfpgoVkCYgDaV+tW30hW/N3wDKD/LPqPISIsNY/aZK0OBZ
0XYRcRRWWIRR6pSnoHDPFKFhR0u/YG8mjn9UutVHqUgG3L0wL/D2vcOlHA/C8odWltH4J/Y4kxc0
vgoSSdRKH6fCANKo2UOgEzUWhnRyH+x6p4hgf2IWFd5T6B+QSQECVJ6C2lvutOJOapsfZTEDup+R
8gsAe289qOgule1xjhmWTFJJpIbWs9PWF/N64+kMMeleyTp3v+1ghdDuufEXBjxHSDgNgrdouuKv
70KM78q7dDsz6+5wP2+iTSSHaXwS7yTDnxxXh0jIfMNrfFBnF5TmM6xEFj+Vm7fHRGV/dXWJB4I7
7RKyyyvnacXKrUhKgOqq+N9q7SyCo6vDVK1EJ5mRkxXW89/eUdEzLBgqCHVZE/tPCde2BsaKmals
9k1DyLNofFnfucaxY9TNDkkuYVO04DpUKDi4ZAA9arCxa7duFssqPiWp/nDSKV9vuGwIkX35lmMF
Ih2fC22WABb/udbaAYkQmMhQhBON0yczsj9AygtPUmR5pKZbx6SZB3k6GNPntqnG3W0VexUw6XGH
lq7qtoxIzmcHCruy9eNcHqb4hQMZzTd3TXVcGxsNeTlXFR49c3u00eA7GitPDt1J7aq/N/z4k9hd
YJWY0Yt6Y+yStNjjz1UGG144asYpNwkBRtU5iRyzx7JvxGLSUmz/SWOw5Ti4NmnKNp/Guw4zK3b3
BRb7V2o8e1DsS0QtVUh0zqzAxEA1iKTns0SfbXte626nAnmBoiJMAVAvhIeFSdbGeQ4CixKDo0J8
RPAsSJfzumSxR2zaHqISxB4Rg44TIE06om52vBMCP7Jg1fx8YFeRoMNqTefl+OWawJxIZEDhb+is
Meir+PAbS0r/x+gBzuEb8ZFaZX3wBk3M9DHWvGsMJCPTuoj8ATP+53/sanJB1TL3oRC0IG5cTVd2
ZF1obhEpSGyeJVd3PSmviN2qCUKbXEdfnHuYgJ1MVitJc09Ks0mnFL3pwI1B7qzPS+s+Sz/yXOXH
+Auj+thZwOUDKJc3t0znDcMtTvIq/49TP9HeryZgmmjCQpletjYdi100ZTSM5Tpg+KxUU5ylsA5p
lenEpT0xkFcYNTY9DFqw++Uw6s22ibvcO/sqGVLOPGgoGr5K8VqXPz9PhuBKgjsYgEC0YSWRzrtJ
71XU+HRf7UeysFmgceX+hAbAQyUEswXjE1/8SB17yIm9wZeyR9oMjqJxPIqCH34rUDzyUkhTdNgl
gVPozVP1lQ2GG1BE3aTIpIn/kI5SivSoTcLFJRP0RLRCMDP2+3Dz11v3UGJObezwOYreeWvwR2Ff
YnqEOCC83qHTV2shCXZAZN2ADCJjcFs2XZuwr8bEHdaYfEKTqDp/RtvDEf1jRfINQH5VJ/J0srXc
UzjnRwUSy8foqveqVHc6Fo/uxrrJXbnCLvOqBCr4xiN5jeSCiKolENekhm0GRB72GPZVFoYUWVS2
9fPfZ2RRnE2fQir92cvyZvEHBTiM19dQH02CiILP2nrcJCAchkc23CWGVSGCwtz9L6Hc9jTLPyAq
I5UmtriGyFezSHyCzE9CU4knZJu8uqnAWfkkzLCZ3i6P002qUxmtCs+OfnA01pZepAKKdpB58IVs
YM+dpjoi4KISGES9BPhfyy5KUYcSVH7awysoDZ9wDWq44tYn3Lcqb/mO15kaiKrAVMMYGfzUyQOF
7Q7YVYc5FsJ2U3gSfF/Ueo+rLeGTWsBDSbXLzJiymaH1QWhJzW9Hsc5T4a1nTqGbP3r4qw3ARrZ6
OqBfywPzZQQ9OTQ/kN848uxWfX5rWBGifTrqgfdbOo+X4aTG3eM5Z5bUjau7/ho/DqtNxJPvNrLz
SfoAH7LfjQwqWUf8h6Yr770deFm8aB20TLX2w6R1oh3kLwBNMZmddfQxJSLByqnQxn/t8iyLo2ST
T6GOnBexY9gmnZx4aZa/R31m+A4aAv9Hf1axtxIyfz2FVLgs5zMb388p7UWWROhkOogYcciksvx1
qsaE7rB1iO3Uu9RwT/ceSofDWAQfYZ7uRSdD1bI9VvPJYwZpxDhFmvEjPFBSey4ddavm38pWTNkb
E3bPOS++bBoiTPpK/e9rf1TfvDcBXEI77kDr8gSQbT8j8QIX3JC78Tgrv5ncDKDd8AUx5//DthQ1
+2c+IKxeVJ5MealHaoCgvkd5PsN25pdJxplwIKoly7XC1DEpWYapVg5HQrFrdHgiEpruTz+mrj3p
y/OHXsHvj45kumO4h+HJbwjCtfSJMF2kDhYE8iH0bYuvxID/irBz6uuKMrdpilrSAmL1XVGxY+Sr
TSoOwPSDic7kl5yfH2QK1tMYqISsuwz+YJdEhrnfv9+v3VF6aJ36eO7auazw/sNMQVRlaNZjlzDl
C7MOkPsP0EyG98pQMhB+/RpMLqIc0Vw3/IFUbSznYIcOnc3k152RkpPHSJBUHFMimrceE7i3msmY
zMNVx/oB3J5KJY8cMSLUvKbk8DywqnTwkmDjKHZwj4p7KTO6PuA59rTUq+56eL4b52n9UBeKnlic
b960z8pv/deeaNBOWn+Vu8eYx+xpNFo0ZxS7IE/CVB7gOU3q46njhe0fj5yMO8CISR2XBWf1wA9+
BYJGr4T5C+d/9azkZ+M894dePaGu1u1SQwWRNcy9tldw8NMToSUZ2Ue3OPzYFIn6G2goexA+Q5Le
FRtbunJtdfobju9bX70XChbVbsfe84evDkrEEOly/OGlg80p8AjPMpjvONmT10o40FBMGdArDYq0
lBwx0Tg2xKi9/M4sGT82iJe4iVvNY7JpKiUKfi9qG2XqL9y5NraJ/qwYkxCIRj61Jja1d12j0FQN
1ACMJJenAZamnLXPOGBoLRbGHCkoOkY20uyrJhZjasA6ekz9GgeQK5AFMpviBzTPbjiUfpQiYSn6
7035w66JudLl+fyHOrmEWQ2izKuERRvD7p4F2CbxS5IMj4+kXXJRhDDcvTxlxqzGUttGWPnu3xTM
ITakCYJ3V2dBSb+LZzeg6jMz91bx0E4bh36mlyeEKmHro0y7e1lWM6QGSm5UqkGHYwBRkjSrmc/s
YhYLx7hB8uPNlbu/54u98w7zE2LnCEOJutCERrAitY91PI3AtsE58wJ3lfL2136W8PMoHnL+9jAV
XuEuu3n8vOYxLRukzfkg/DOUloLOxuI8NV7wzpDi4QXJe0UG9CsKqITs04r2Kk++r7vhEWXqP9pj
MkPKxlb8f9xuQn/kIpqqV+E79MXZUip9obRuvKzObIRv0bDVmxwiQP+sHvMuFxMhm3ZShQMlXOdL
e1gJ/LOEPxHGH7xxKSS+v/I+u1keb1db77oAI03KyDKf433ubI1H2148hq6T1MawXGzEgJ+86vTM
LB4n5C/+YmHB36nFRZEY2d6cQ3TMSTZq9EtT7dazeEMjwEfuh+zgKt6/9+HPZSUCNb2WNIDNYgx5
ziyV42/eDfylgPp9NVDUzn/W2ZVwmbweXN7U8UiCFhKXsbeDkFOzQ8YCPyxivH5WTXNckZgyFDGW
MsQyySs6NyTzDmmywI5JruP5I9vD+2pszoNn4KGL4wwEoP/puwN+DkIUKyckbBKSZzSBqAeq64hE
g6LmyGPJSJQJCw0BBWAX4pFDL8sLKzOhXi0RwP9smkdy1JU+J5VeQfuoLgH4EpKArLVpwYKcT9Jc
qfUxxykhWLOtMbElY1uV8mFQcV3VWeYPC1aa1lGTSDs0d5coCoWbK5rJRf5/sLfC55oqe6VxrzgH
gAl87oqCtxHHwgIbTeHurCXv2gyTsHawNzTDSwxstEe+FSeoArOTl6yDLQmrX+gTa5rYmSoANyOz
YES/qFqZaVqw3dZKQ1aoWXwcQofWVoLMraTU+YTvPMwXXyK94nZRUKi9jmCbj65M+I+c8MXruPbk
VtFPbsJKiN+XvIACtDfVWVS9J4Ri6eqdrI3cq2vMPNiY8B2LCiCOZHQTXQTPKimAQQVF9sLFjc1t
/0YnAvcf16HacnwwQ1BpaH/Nk3w9/AJMJ7fDLNNtxc7IF+u598QxXrVgl62w0tVxZc9oOZX/pXqA
zGIn3f/dlWO3uswHeVcTU7eNkUVbSRtZPaD55Ma/hx7JHMjAVRA7OHGUDN80YF3xXgLxvm5KgabI
/a8mgSZqXKcAOzqLYWLatp2Jggiqb6LWcppmy0/xLf3dE0O3hKnx1EnZ8i1QwY7H3u4bDhfMHW3X
KgaHVwSXCz5QizdMdrzL8+NbZk6jGhQaC+o8h29GDJlUV4H2ZG7snSDyFdlBk8q8sqHVwDLCTuhQ
zZ7JCnFUoNiUZuwLemU/STCia4uQ44recchwfbD6JpbQbXsswpdX6eTwSDeapUbNv13gvSPsqoPP
ya9DCoPbha3me/UAUTjnGP7k1IXGZdspDT+DnQ9TnyqAm/uBbF10j8acZCIKewnyLFGY1SBn/yJw
WoMescvM6QJKf58kvizV5/0BiO4tUu/nUXsmpuDZ45iN4i89jOW2Vhsv6z7OkladOLu7rSHS5o3h
K5cAjcyC+jg4KIZ7SX3hwnp9GvtvKEAMLfgTX6EUrUoS75NydvY7dZJgIwxALM+XR2WAM5GkZA4f
2tZ/7BrBTPehNkNMmyKsGq8NwoHvqsXN2Tj69PNNA5DHw3FefaTetrgbVjB+3WSTG86ymxpSEqek
Cz8dbJZUgwlX3IKQAUZNZD9jqZkf4oxrzE5IseE189Vqgd8smI5TggMiRkzIn26yFhWGHHACCyss
1Om5ULkYSAsmKMW9ZZduOslkjResY7w3Wf88chGhMp+Eu+sx7sCQZWWl/i0IMOEiij0bbL15qC6Q
bQ+MKLnObU4jiY4LKK5EzCm1x6Oc9bEkkoKHP5utMF30o7Vw79limm7GYacFqa8PFi+B8wsFzJXh
tfC0SmdIASVMHCJjhaXuudjFmpIovYYV4CxIsx4adfH696ApqrOXCp4esgsMwJzt5lo7duVNXCpM
stRZOmVp5NLd9DRHwCWycPbKu4zvJc75WtdWk6zxcEqu6qWs8bx6Eh2j/44mLc9tCikYH7bKOD+k
zTkQC4O7YDhFc84uAq46AQvRRMs/rD7qiQ+erZ+WXMA9cbivpfNb6cAt26JjvyVrf6gW8ZPhOS64
Ldsywvietdp2RBROEzRM5NpeziBRuuJwBTjVRp3mfIYS3GH/3+J8vu3+gMqy55itKwvRGyRX7VwZ
/YUFeI44UMAnrMdIoljRjuBt+yj1EOUgcifnjfjUCK9RHlGG1xnz2gyIR1HPByAniq7G+WiC5OY9
3uA69wZfA4awXjtRl+su20pHqfSdTY43pOc/oHfi7apG9emv0D2VRed1g8oW/f2fhiiHb0tHFQ3i
AvU4vU20SnawuQ01i5H/jShBEiH/yl1U5IuaB0KfLMxMkmNltQ4qbMGORqO7fGzL/Q1Zoql+4yLc
rbRpmH3OJA/po9WdyHdPc9mH/gO5yjNHN4VS6/OKEyPAOYO0L1+JsKyNf/cyutRcaUXVtVoAyYSv
FoQ+Y92CuRTtG5TLdo41IjU/qWckrHuzIrdxtNxGRFYh3zq177JORiGED4icddeChtcL3OInZRcY
ta5GvoQuiNvUZReNrfRSybAu8CcCZsvJNN+EXNBKPrOoOMmqlbCbWQAyWWfryg5QNC85UkY5Pa7d
LXJ3SDW8GQY/lbdrs7QCwmmwYVeMz2MJdpo5yUiNvwSjkvLAOxTrt/ArXo2f1Nz3ix8PjSlcedzL
RWbDiIoP8/ud7mdiAb7mV/0IOIb+1hESb7Ln5zp8X10ej+JNCX1YxKrs2VgwMmoLrN+lIRT008Hp
Ph2GMyEf0M2xdqvKN2jdNQgUuj6tmWWhL4Cm3lJh6qcwq7X5SZYIhvV/ftVZf6Npor/JFLpJfHJ+
G3XN/1/fbvCFI0jyUx9c0RIXGwYYXf1Lo7LGazGihoaIWe5lnm/tzD2Pa67WGWi/vMk3evrjMLLT
oVoGws7nqIJlrjwsKpWfFOhmOa1yGex6Y4YTKZstoqFSBek1G/xcIaXs1G94htU0sshsNIp9z8Uf
JRt8ImdQJ4SpjEJMb9vUb/6hQE4hHvLAl/0DJJ4DCrQ6H7JE+yC03soFBK2GDgan6lB2XaAMNcKw
YEquKNEShbYXmhWDz6Nem2PaI1N5NlKk6cp9JkSh59buLtBw74cg3+tpGQsG+k9m8lwsB9WJpAuC
Q9o3gEaKkrYtMVJf1FTuDEULQPcMJY6SShWKiYvI2xyd5CyFv2ZNYCHQ6aaakA56VIYKBnkbp8VB
RyUhPEfJrr6NRk0cJwYomDGSKm4RvBUgHTqsF8Dh98ErCAW5poFPkO0JbOib95cYAZGLRsO++yN7
sckzfCt415ng4Frp7x9XRKYECSr+2tD+amrthA6TajipbxhWYKGAvAAGsUmwPTUUAn69TyY289vw
rRqVYjzznZqFKuv9/EbNgAfNdTn5ziiNmxOVS+I1T+mNzdmuhQtnsPk8BXdXkF3v/OSj+LM3JgJm
LF7MUBG3joOL12Cf3xGxPEsRt+NeC8vGaJzwHF72i4mSzAgm1yuZJBpEzH9mSYRFCFhfKj/qwyxD
9SzliaE8QzEgaAaetwVv3R/t4nEX2QkGU5ddX+nod5OAfzj9d2Q2E1S2FVmeJ+if2uORTMCf+yhr
fwv//n0ZsrpUBmYi4Jcj5weYSCdgJqmBTl+3LSRWteYdio1ODvWg+dqcS1XfL2tZjmfqKW24GpLb
uRZysuvzOY1QZ6fn4VZhe47rcMDbK6hBL3R4O6eV6XLaCqrfQkCr2JhT7EpkjoYubpcVpWMu1bGP
m4lKOYMw2LKABTD4LuyuZXDWxMX52fW43B6ICPei3Bdwar1g5ivScQPZfyiKuqv4jl5OMd1B29VA
laWeunvV0FRp8JyzxiV/wkIhFZBnEdFvD/SE6u7nl/eaRd9+tf3IPzs2dC8pip9dlwkDxmyYVgKi
Y2U/LpqyJWfgJKRfQV5/Cvh5awWI+MCWqKBcNpbAZ4+yW3v3IU/lUDe8YHLVeq/XiIMdgoEIGfpF
ceg9rTQH27vw68Cr1hHqWXl3pOgM5fdbIljM2Z6FwnwRPKBrlr8eML80dCLDBWMw8QYB+dX28Ppw
lr5d4xqUfFWaWEWBm5EqEtmsaOyCmnzz4g7xAwKwfcH8TcT5SyEXKltNVAvHkNlCpYsk7vO+s3Xq
XGv5NLyNtC+3my7H/22hzJLU85Ei4CsIk1hr/JQ4ZlhgIP9xMO364BHXAvWYaENSJnmGoucs+zkN
TQmQ9hxo1gY8Mk16S3Z3vFibpmMMvSMeEYAtkMGvMEdOw/C/wKrngFGS6ZxzD/0XNDzfQrzYYbCZ
w2t1P61SSZp2Ha3iZ6i+M65MX13qGPnu9+3s79AWuQ00XAwGpusBdXA8pGSn+xsHIZiy73XH1UmH
F02lkb+6wUuXWjkgALJhA3btlvzJaSnZgdAvIUAtd+71uJiEDXrDD/U3IuLPEcd04fXdHS7FPfOR
5AHaYbd3wt/7iPDBuVJ7tjizbhR9Te8/ylaFVOtHxYx1laCVZnOPSTBiJRXfCgke4AAmkrHFoJEQ
pJtdZEghs5kr0mpYIFCbH61ZyeEf9PgevuqSUHdERG5txe+Hrqi8RVGQ4llAHVVecpmlyRm29Qk8
UdhLGc3ki6zAZbpPpa9oxHZoPD68NlTWJUjbIqVpyRyATzAvxuP0VvKE1S23FTxnRCvPzRZxXonB
X1eY2ep4gZsCnb0LJDR/btmJ15I2M+pcX9wg06GNCz2fgc7Y2pDYb9PfLFBfgcVTtrb8ZP3lUnEy
MMmecbRs8NdOSpOcqXF/FX02OOf3Qp38RF31QyxdhWYSdTUK08t5+eFi8GjvK15L2Yc5JmOKUFNb
SvijxMg3aqmLixpQVk3S726sktjQR+Y/+pHc8cqTjKo9DefUBUvEC/mvZVmzXlFJVO0DEXmHXJ3A
YbpqVxLrdNTWVg7d0KmqhzJh5X3GbsxqA/dKpbTMRZboKjPxmkuPcWlxZgcMiUT5hJlLdz7uDflQ
eOLO3kFN6WK36pDNXPwoidqIH93iKxRDk8f0eADR31SNuNHRiEs9tOTX/FxJ4yvIuGb6LRg62lMd
rhTsFxV+zAO/gOUgYS19E7k24WmsXh+rbmfERrZsSt5nPYub0NUwvR77GTOfCPy0kw7yRIP433w7
rRw/hhCp7XmICLxyT6fGlMbCsP7WoUpGBY5XqTlShv81LJBCVAW8n/ue92mhuVRPnDO03oux5+V1
l/aol/H3QplH7XfCt+/tzekJfuxj0QOU6HKNMLAKVFTAmahZLPXJPi91H5D7FDfNjNFXFs28lbK0
sv2zcO2LaEBMfmiiREOAHN1aI8ToQwsZt5rOpoPoarz1FjWXHa5vkrvvCqxdMHT45FaCt62u3p1T
sgoadEfp8dQTZM4TGvzHNTAoSCMLg1t/r39JcVGdOFjv7Ez+YAVwsdYPeIYaQJfXqCH0TFx9eag+
PNKhK/ZscYDRxzV7Hkv/wLNtIxsFfFQAhERlb5BCqRvppgJNuhfKOxFn3GTkiXFACKMoWgzwlO1X
Lr7RsLXhN69Ho/2KgeK+QvxGhBjZRYAiZ2vAn4tz9wn8MPU0jbz73u58jgY0MKIWi8okKYh4Wqbv
k6ulhzZpD21i9s4IJ1FZvpKNnYjDIdLM8qNXP6ghueSeNnt4AafzHYwFd/ZWiSetNbEnu5hsNimK
udrhposn+ltONQyzCAgKobxFpyoJfisVPk3Ch3hNWz3LCIEpJnsgdErBSlbyF/xjBc4amQfK2E1b
srCdHfU2s8gbGs5F1A8f78QrVbIv5vSD2f/Kft+Clm6myK1e8ILY0nH5FVu4kHA/SPQqmXYPUDn6
m+fp6n31ABVg/u7lry2+cqbpqoxH5TnddtvJ7HHj1vyw76KmIZkhqwaSrsKM6NmAPq3eREF0TdG7
szqY+Te/ZGsogzBpwkLYmz2ahewOCLnSKgh9NdY7o7SoKyldCNRjvWluEW4BRfgtXCJq5EPFQqMn
QHjcqgQy6REsuRgfZT8Jtj42I9CZQtFaudhKOULrk4daaS4/QMlQLWrg5gB8oYC1u6p1xXl84FFZ
O8LzD3uQzwR2XXgZVy/+WSkG0ni79mhmCEbL+I3y95ivxYn6oBMu+Ye4ihL8YiBEjrlGL6xYV0LI
e8hxCVEx+wImehUcJ87biE/KPGp9IbzCs97eWzfqsP4w4aqGj3pjyhq9CR4pKc+R6XfbUE2DTm4g
Hf5ug0Pc9duYFz06U6JikIr+/xSs/IKjrzsHcdQzASj6Yeav99QDhRCcf7dSAjSaw7iWaDu+oDwM
BwqXr3AZI1XYBdLmdi7heExhCq5EV/ROOC0lrLbmAUOLxw/e0vv5KM4++yU8xw3IcPvLOuixCV0N
Y1f7TMvP+9fe/M25y0fMfTOd9Yf9h6mmBd0BsuhBC0cNU192Ua9zy4Nl4BrVUzBXinQL5Fev2QCs
Rx9Fjzjt2vy3wQxidp79oW/5z5g/z/x69SriA/JvlAlQKS5uycpmmNr7FLL8z/pGSXPafiKNnnk6
OvCS8YBRccNyqb8KQiq+8ZCVfCEUGRygs1kYnZN+N/Gby46nvJZXfFjIGgPkHH++ycAeAHiMdq6t
AjhR30k607NQVS70c4IebQslmD9h/MRoJbnFccjZjg7HS9mt+glU9eu/7bC+wTPx9YmfDOCCmQca
5cp40MUKShZ+dllGEv2KF5B10scLhMwZahyG6YeD0+5E7MG7u6/M5LZ/3dAl2mfFL8RL14hAKCKX
SLC9dwSG6xubZzvoz0CDB7py+G0A9Ji0C3WxTvOajJq50T3PZv9y5F7Kg/mULXLg4SMaUz6fF9AB
O58nq9T/aalalC8y43HR9VrQPwML3MM9O4rHU4awTtApqh22nKUz5QXr3G7e839bkdhUVrjEHdVR
cSJAMeZ8RZw5R8rYudNNehLv6C+JsndDGFZyxbLGZn97Wv7N7nxRrzRfe/U9DH+LwRrVDcVKa/b7
XVAp38N7BGOMAkcJwBeUuxcIpvYE4nadHyApq9r8/4hzO8WhR1vec7uHoryDvRKeNNgw4pjGD0N5
duXuPe24rQO8JIvV9HeptAZRi/16NLwF80xv0deA1n518ZmKpqV46qAknwUyk7hrJ58v7CPTodtU
X9FTMhz5S0ZtkF1IjclKPMpawy6J8TQOakBw8dZI8ATxeHTo5kzfmEzX4FXf9CJ3v+zQ5ffZxN2U
6ghJsOqeUOntJvYifILVOivTBhlWEkguUPcN6RPhbbLG7Kn3z5QB5ZzGFtANLYVxum+9+wZCdbEZ
0j6fmloNq8dURJ/6lkeyQ0Z6xlVtLTGXldmYKts2dwHXjtSiDeAX3xAgH4o8tE+RmmVy3Ugr+knW
MWtQQrXfkFXwYBH7bNqAMYy8DBehOvtOt6mBMncSzQVg1Jq6PJ7u82QV7AUWXiULVvrA6kirTWEH
UbgWk6Av9CDDlb7Fje6kK+xZARmZPhqcbJKsHHLDTUdXbN8C+bZuf8XhX0k1xhQc3XYvB0BwM9eJ
QWRw2P4Ph+psR14YXREPWYIXOcY6/gpILG7bsHPI+CRk4idbGPeUJhXdQuteKRxQXR8zzSAjpl9p
EiHwCQTQYCajICJS8qpQXtMFVfBhl0znaweyqjW7OIJNS+1NQwPFBxjYNX/3frNHmqO1nMMzJNHH
MKVSrZmR6rbaNq+9l+BlrfAmHhOdLfBPXPcC1a+mp5MqUbbp7fInG3mBVKPW9ByyWv9v5u4xv129
OgkvevudeJrYKC55nkvpPtY4y+jYe96kXZVv0V/KS08z8Bh56gk+wNUxDifjLxuVK2NMKoOx5pCp
il2WPsJWo/veMzoqmP00CQbsLAGPS9hsnTrEO7OFcRwQNEP2A4DhVf/it+CIDCAGaAYrpTTUeuFl
liQFv5qDxAHyStyG2kHL1znzZBKy6jU+IOfKBCUM04auyl5sRhMX6fUcOfRgPn3V+V+aEUuNF+y3
BaqlJcD9PQcTc7HXDk2c8m1qgzc6jYc10KACJnFFP0s+xk7T/f2IYMYF5GS+j0HOstMNWck7ChbW
cPDbWk3sI2Xvpbz6kZBVA2yHWk3/zfXHnhXcqcS9uMesO7rlp22f3VZ4W0X+7UcdW7U2KUeWqVon
jCCN+6e+sfpQEZlGkmE15Sr0D1/IbdmuQAtGi+Qvl2NybvbkKwayCCcrQHmW3qyhyAYcTyP0B76v
dsbeJ436LSawU6D9vh0p91HQIUJWumjKrDjbQDh3LGy0uJIKKcyFzUriMoAkxV7qe8NSM5yWOfPK
65wL2rxD17stLj9UeqhBslHyZrbdvdnIIgDDUe3sxlgkXnjixTMvrmc/TYNHyh3/ZSJ3lPqTjVXG
s1Eg+Yf0AjYOL3hvNfnlRBkRRgjWoniOzisM+TNH/Gp2VFvSx3+FagUR3LRwZqd+88FrF9Av3Vu9
7pZYcN8UQk62kXxz2o2P0q0GJjGaT8GG+1j1T/1JPCV7T3KA/JQRjptVzcVPQktj2hN0UrinoFfO
DYjeGZnSUnnyU/eyC7IHBGNqneEu2L42y/hzJQiquGUDolS2uUIm0mIKTjoM7NYBRBV/RJdpPuCZ
jtEXHpgmGnwWN5uTIebNQF9eMzfegAVEhKh/D/TOAlFePwmnwPZ6O8sKEXE/6oicU/IWu7oC7dqj
HQmUdOgjRAhhFkVVVntaGdmsuKbKA/vBSbYKr6lQ6MaSfgfkh2tvKmtQKDvbvPvdcjmU0TefE0SH
IwpFubGB4dAQtUjbFgBPcYdLZOk7KdeVNgt3U70RXs9k973LgeY6yczjmpLdrIKYauKWH0VGqraX
Bv7QaozHoQk4MuqfD8anXkGLTN+DyAwgj6eFE5qrpHmR5Rfn5P5Pin+sEdp3yfLyo/ZDHJhoexnc
ISuLCdoSNI2zyvVsv2Y/la/aGTf8tgGf0HoBmwLMgYmtUE/iU3Pr1nDRxQAkpWQsHISIiGNLM6Tj
mcK+ouskiC2R44IvGPNkneM7KtctowJypLPDhchDkfymjptQODmoS++O/VzYVsIsvWIRhQpRt+Hr
4SbJvYzGYyJ+MDVFgJ+iS2pieZ+/Fy9QGSR9nrb+9XlkBwtX7ZqbDMCMqNGtsHk3kvsQr2iroFVU
zgiv3KfYIhsKpteKSBTb3G0irqSbNQfX3azH5QUU6/MSWhVFYOAy8gh8kSLYi3Ej/sfSQAsAmAD5
GcD4inAwhx6MCPzxWEikk2uJCEl/BKAAeqsq1Y+dnjz+cOGwxse+/AzoNvROGxiBpJRKwwrPxAwM
zcr/5UnqOA4aa+ijU0XMg6/ABfSYSOR5ZVWH4Nx6xfJ+tHugAT0ilp3ih85OD6A2cGDg3H9w0vDB
zeVjLAd9Q4FaFRdNbZAB+aQI5fHKNVmDo7g0Z1xJl5eofHBZ7KUas67v3Lal9USy+l1MSL6nznIt
UZ4KrCimAIPfiBaCI0JFfgS0Q6aENsV5zXpK86oxlYofQjI1T4+n4u/K9oXXT36Ln0W+4j1Y/SET
wdS960yvHoB5Fn1wEVDHTc5z1x1/cYWRjJ0XzTdRxnP8jMM+Yi3Fb6CenGiR+AfGAkEg94FJWv5U
QYXgft70kTQ+WOhmIXDPzd5cKB1WON++tyraLrE3rrqxkXmiBfrbyhj4DCGSIdl1+KfwoARqfUAv
dIsNtSsxDHvrsSETM8wTtdwV4vUR4V2QQ9afOqXzN3lI7piz1mJ/ow07FnSuvMzsHrBype8MKMDV
FVaQVUOrmtRnjPWrXj84/PbBMctHTB1jABIkYUSVlFwJRTJjDSR2kVGnBQZjo2iVqGHz2ml+ELVm
drj8th9m+fKqlKVGRWcwx5D2xQpbvQdL35q3ynaUUBwfDHZlpuQvxPSYUrc8g+hAQJAjU90gg7P8
1BC5FDYh9OvzbZqLneshvx7g+hMQEBdGyopARXZeH3jM/Ni9HmUsIsgtj0C/YOlfhEF5g48QehrL
SIQbDvjSRz3KluY6GTLdxM1JybmDyQjC1HxX3QO+IeyJbxhBs5yC5kLPlI5fYtbAQLJqOdFDKTCX
ulwJvVoeL5m4Un2mECGHCCsExtt5IW8oWElEy3PRtQ+dBVTzCG/9HwK5qVkfdxjlfPjuDs4EXKWH
3hE6of/n/sRh5MSfOWnf8nbWW+BpzDPUl7T7/9opDeaQyRrFB92issYMNBrsHosBSn0KHGr13vuD
JPFnBBHgqz125YW2C16qZ6fvQBHOt/GqC4plfLBqdXTTEIVMLF/EJf1lfONCgzDMyoF5JjF85rVP
N5CNkYzhzAou29i2F/MImswxP7/w0s6lwPKfjdq2sM5dv/jwZhB9jyAaaorLqt68U3kpIui1H8QJ
O88GTNBveY9xkm48UMNfa6WKvPoJdzgDPtIvQNilzWJ3ysK044LIPQ16j1GNj2Qhcz747OWdxYYJ
AQbzYMQskqFogUYw6rEtPcZFh/TXU4+yRHf2cvaTHY7TbZvQtcWnDIL6FMCQR/CBCMn5O2Phj8vB
RywoZsffPq4jZTXNWBVujY1w9YWQ3anJdrGDqhImYt7957ieHICagUW4BiKE+D3Nb1j+1oJpMMvM
bbd3vrqkMVw2OZcMxhlGo4XUWZedViPnJRLjv43rZMRW/C77ugoBLfCJqonMlXDAFyfE08pk3Lgc
Kwui88CtBS4yf68vfIZiLYCfmnp3cNciUOIJn9WlKm8L+068fxcQWY/F3/bVgNYDqPYuBeqeQc02
9SbXAB4+E+kDq6bVD8KTd9HjOInKhnOgrL8kAU8BPz3hKb9wEYMNPxPJO081wGGY2fKKoQ3j5dzV
+zSjFCmBAv5WAIfZ8Gk6jHXvpMKw120DxgO7J9/zITmpNtfBOF511zdUkahag7Kr0Qe69JEE9m4r
gtdmnSYXOUdvNlBnIZXIdMs2UOD1MI6LddrClJdqJXWUkNJ9SMtRHOFxmTOgj3smA8o6TlX5e8rx
0db80t1Bw/ZUzLdrJ0AvKlL6DMBXPgxLLBi5oodokYXlgePkMgjEQNS2VfrBC9dgZaVgQx3badoF
BTdYRJMoDzOSW19i1Px5pEjjK72XOvujV6TW6+R4g/IyMI1oUcKjfEjKZhZaFoODGWl7byFiBr6s
2u9ic0se2iaWld24wJ5OcjUPFJunpzw0otJ1W1agkoQXOiY3iUSxRknYeJ2J6/knrZCo6FgukF41
ZYiCy4EjTYKG0gOF1+mD5wnQ9CY4+DQaI6Rld3MhI3Csh585tgSgyL9+elOzeYPqSKnYBz0e3jzh
F0EP2QZZ7n/6qz3LqsJkUkTyYYZk4Srji0LL9W7BAlRuiY7nfQL+a2Nx3AtT4XmOdUJ0ThBDJuIl
DFoQ7LrGI5AqEe+2iGBu77PGjje93Op4pCyRW6pknH8WaxLZ7Eb3jhm44S8ehPxvCYLfkd/K9DT+
45sgHUgfK/C8Ee2H60tUK/vFdQrYzKf/T5ABhQrnAILXAHM7sw0dIB9dFqefho14tv4o5ZI4eC3t
IGvqByMspIuGB0mT+0zzKhFyolOs9WMBFkDdcpCA1Kyl3zSl71mPMc0Wux/5CRW8Bq85L53O7CZi
tfWoIDxl1xaQHzyfdncJnBSao2a2h8vdTHmG0yNzgvgWPo91sME+6ULLdYIn1104Omb2P8xR882z
qw7ljuJm0UE+5k07Ur08gEvMTZPiJlF7DYFN5zOB39XxpvOWlZVxMh2Wc8xstpBce0/QGL07qtbC
z+TRmS76zKH9HEqXQ2Oucj4Um9Ymfp7zzcGw59QrSCgZC3RKnthj/VekWJLz3ip4sRU9rO/oD9hy
Qt2pkOC9ycn4+1NkfWMgABkQKWR64Oz8Xf8rWBz6a4nm4TSIJ9iRgvvWnpzjMMQFlAFCaq0R/I0c
Y/PZjQye4/rtLlMACqqQurmJM23IDA379dGnIZwS2cuQ9d4Mn0CmZZ2fckWfG6s5KlQLdNvmx3lv
iFBWJrV/bOw8QtD5p2qNQnQRWMtsziulX8fNcNvs7Uz3ao+KtdxGvvkdXfx1n6tbU59PvQmERodR
LUwtWksKNYFvTY0y6DhUsgL+Z1t1gH1kE8uSzQI71q3VMhgc3k6+T6K73LcjQSzxN5iAP9M5Msxt
g/NJnNsvQhc1IOyzKoIwMFCv+0ZdX+iMPgCc+AvlCK2dH+LrmDtCex7ylOkPxTz9ySp5leCA3Nge
E0pOhzh5Am3eKNyMvsbNnNP28kRxuv6/hFG3d26gb+aWKdwhrqrtd2dJtOX+FfzlW5ePnC6Au+T0
PLCMVghjo7OadX18H+w+2zk2omMFTEtLEBLKjZHX7ZIBWjJ6OrOos7hwPUYNmzSyJ6cfdn4/hpAm
oWiERVj9LsN2c7tU34QX2IEILToxkrlzg/ubTraNEqFmcAwjyrdXG/90v80+HvHwQqItr+m7FMXx
x0CYrWFYeMF3EeHGEB2cijttlpdczH/0W2RAK3acN9WT6OOWtfaxVE0xnKaUv6a1ZcNpNez70Fzg
IvLw2xXl3s6DAd+PyvfFKSa8b+us3Pu2c1YK0eWEZ4Dpu/4tbBPyRX0G7sc3DraP0IW96Ja3hLDy
pIz8zT1HEgltLMWkQP5Bi8bSUdFhK+uh4lbrbKzNavKuA6Nv4sDmzokF1hEv3SoHX8jg7PUWHISI
mm5E5XpPr8zICfjvC1iJScqfUXMaLo+e0hFhXSAGA7oZDnt2PncX4qge2yjEcOFP7F8B3wTNXKV0
9/xdwz5s1QQTgyfzgtl6zLl5wRL26nl10i6L7cxa2nld/o6nIWi9pZa2EJVkQN83OgaA/05QMU22
iIs16WRz0Xj8t+x6IAW6ovC+mQ2Njk8cfUr/aTOhn+MuFDD4GEQV5w1R+6FBD25QqEk0JxhvHtL9
RM6SVgtwbv8+pSwK2ndci/u5zOPM8gkWa4WngWXPRHcQpt3/kKTvpdT4yo35Rsl7CtZt5RbHN9aV
yqMGwM7ymx8lRJhWF3iM3N89X5amiDw1uL+HlsKIVFgAirwzL1+2uGEPDYQ/SamEmn1LWbC27Che
K9Eq35VfQNQKR8S9kbvub7BfkCtuwW0THvKouUojHD2KLUbmp4yTSD4tbL18MH+PHnzeA5R2ncR6
DuTpeNTYwe6bDlLg3iN3GBnNEHEG75Zg1nZyldhyHu7WlF9CiSFYHqcJajxfEuMResg4UtT0sAq2
Pm6XeeszUXA5D0ADnwBvvYYxRWWLE4tVzcdz8aaj0FFasgxyCmSNcV+/hEiHNtjdJsfqs2/a1RfQ
BafrLiwm8GMQsXeZlCN/fs7uvolV/+PGkMxyrw2+yROsU/snusx1aBNK0oSRgIZWspMoOw4yrbaH
O6/lpCfl1XhwruOTocdfNKdU/ftkJXEM2G1rIInvAoO6mdZbCiyDhSyjK9o1em6vVBQMXMMhNtQh
BA3EtErslvDH/99DEEs1bQP9RbXvv4pkyZ7d9ywugYYMbwF6rxaZOwGtnLIvGWLpN2Q1oiPTHwWS
r2stzBCqGn/wILEFqx+x5PRRq6Cl7i1d1u/CnNqxDDfsiNLP4ZcfE3xYDBObHpfY847B/clCL6ER
38sYmUuV7hsLRUu9ko/I8nyQHUojO5s8iqEzZtWtgtZsZUua+K+8669h/86Xp5ZkrloL0jDLB4Ac
7UFtRvfxBznEsVyBq6n8eKr1PWvJkoD/kLuHttmwo2MAfxdXx7c0oPKiEOLjvYB94OEeWxkYpwLs
fFvbj4y62SfH05thMIeoj0dBhvcrPWP8xIQYzPjJYdcNT8j+hO7k+qvlwvHO5pCP/XaxBFhfndI2
3M4YWACecFoqmIfukBscKyrMeWyeIXe5RqpKFRyDsZl0xXg3xC3KolmZpcuBeYmQMdJmWUI/pCvR
XL8DVwV1qthti5ntlOeHr5PTpAggHcE23d2BZraj7LPxqDkrwWR9t9GeMSkyK6ncw0NAOuAoPMMK
Toh9ti/LBpf54z3kckoW51ZxwKpdsdKnoIEtpSknJqnIar+B8nb2D6fsdJfh0V/4x4OWrwSD24Vw
620Q0m0Al7gQQ6WsU714FrIb7f2voBrSrDKv7Wh4tYgHnAk9OQLmvyq4sTMsyMPPcahGRNPOL/Yh
xE1574XhRNBQPQDSFOgy1dKCtBX5mHxxiJGzEJ36T6GgTwJGYZOKZGzqs6C6JUsIKR966x+sbclD
BoBrPLK7k8Xp5pik2p16VKQj+4LTvkitlF4el6VA4OlOzWGJEUIZJI2QA8bGCC5FDK7HYNv3DRC6
u/eqrKEG+0s4+WFrG7JJ8UG9fnhQJ2D1yX/L8UUlt3r4Z9FwdPuweuRc6jhTIbnh0TwX8VvqYGLf
B13x2GsfUYtgvmOeV8inQLggWZXryBFs7K7/D/OPemmLa7ZiX8ABvEnUtvMpDqt7Y80F7rMQCKfn
B+WmQSnAkAa7n3BGaf5nl39mXZZxhx1rND+z1kXt8DM8LOQ1/OvOIX36/lgwut8r01Ues3Eap38R
w4hsWFwGMT6HzIiynhCXyWKRvJTRcGUEy32ST0hhCsbm+kbxzGYwn73zsht486yxMCDYPfScow4w
lVKaL46Xjaei9Ax1Y+YsYomp5wll8DjeARV9MtawOa9cZA51ro83WAa2st6AQMrLqEc93GEr8t0V
LTQORCXCFcLluqEm3WItN5ilBEzTdTezYqad9m81AeMJLRfoKcVBc7vBuTL3WAVEPWZbb/ZZnwVC
HFCO3xOOHruI55wWWLEPRRls4csPoL9NuEXxJFCkfPDGvTNaTLWYqCH0MLhYk48sMW1SpbdGzlvA
opULaLxGOCuAb61mgly/jNPTY0wX9zn2lCTSJnZF4cybXDIVXipy/iumETcAHP1DUPW5dHLriP+B
cQWf72IAleKDrnjP8udGJ4HbV6iPuFW4zhnGNKHt0xYk1b9kJ/O8DMy73x4eH1k1j5M6ADiem5AS
K/4k/h4UzcjO6P8+pI0hmpvqw/4iuX3jB941O/7Yxb7ZAv+FeCVHVq+STJM6qtb+9SaPRz/VGvN7
BdoAM4zPIWfNcOgPeXfpUQqZae/TD609c8JVBUJjlL0HrPSdFJ6xAP+LYRg2j7pBJe86DBUnzx7+
oDK4VFMcSgXqbgSA2guJMhZEx5nsoEXuXxo6tblfQTZq2l7Zid2ELQ0IiqgQc2/JPIRjGawqxm7r
DLBN0ukHXN8+HlQ4HkUvaO9SX4PMJqefEcCAb1k6pnMY6JRDijUlKBp69/tpPTQfeyuJmeXVGsvW
NGXW3o8kHMrQvZjTi1N+Y/iRBlbmo9lkli/bPyZ0qhgplE5GzvyjtAsHITETuru/BlS/qMJl18E4
+X46RVDVq8dmZqAE3SpVAhXdeDfdGgHaF5dC6DIADNJBRRT7ocTYzKJ+qFOJs9zYMDid/ycnzzPH
1MOxosHH0eskhrtV91zr8DvE80Bf9Ryiu3fJ003eo3WLVIzntHOUvXk+5bDYLqHLTW4JgdMfq0e9
jlYctTNF5JeyRi8aFaAo2ueYxJPDkh1tdut1hvQd2zKYqCUp9LXtVyK9jHnnWr8rvn47eQn+G8Ff
Ff0TD3dVUN6mIhx740j36shkET2tkl0PFPJSHNeoOzftggk5Hsd4b/zUPn+v8ugpnPFLgSoTvMJW
UvtSIPQAvgJtmz55loUAn+d89Plbau9TI744cdnilibNFiTkFcwufmzePSB0tSyjKRJ0yF0lQdKt
XsozUaf9wKXsoGDGAyensqg1lfbRDVhNGtMQR1TBY3mqjbUZ1q+zsoxEEtJOIg+TM/wRQum3vWBs
jk/fVlieSfuEIeTceG7llFRmepcirDXJ8b6gsyPspSn6ZPyLL2IdimjZOuoEeNgZ3mmmNq5zmLwa
AeQqDULQXpalEt5V+7HI3EziVbwgqRGkuYDBTHexJjeEt3YbV+W6SEbNKJbzaKdAfmUcP9L/n2Q5
2BDZCC6BHeaylEdb0G8NC0z4hEbQOqW0VpzqXf2hpHUdUMoAANB/pqLh/VrGZtNJ5PiWpGyMs5lU
TRkYlQhPJH0f1Niq7Qoc6Ycc+9U8/lGTSS2TV7SMLOk6ZB+M5qK4KeQSDjlssFiqFNsZY0JfGRoU
uDXYTNrbNdJC891zTdpJGiGQY/wDC2NHTw3/9WBqK9yIov5MO5fBeXcKaLHRInpMiTC+FIe3spkR
HFnTk6IW1127PZJxbc6HPsFe4cSODU9ur7d7ER3wYmsiR84TFgmB9jg5d/7DhtkGU/H6VkO7WqSu
/PkTqVLBWxQvzfmn7wMuTYxWwTHladZGE22+Bf95xONEciBsvS5bI+p4NPpY5fIWSUY2hltEj0Ai
6Y7PcouS+xqnfvqciPRNQqxxpPB2b972Whk+smstEdm0AlDTovldEzb9hRge0PYDfPnFuNnJrzH8
ohLAcGQIDzXZy5B8DH7qwGDj3NVfNl1VQw+IoPKEs4wlx9ecLTF9AzOlyoluuHOdY2QppV/E68ly
gBsRXBtK3xUhN91vaBYjDyTEbejL7FgMMFKir+g9Z+pE58q8PjPGC2+VPeY4owuilkKOit36H2NI
LEHwVLgI2fagVYKWUDBzOrr3L2Aw6pLJwLY/44rmHMJofScqpboXDD7x31sahay9cfdLRJb8NnCh
bpJ0FylSOQNvQXs6HiJ7dQN/OTTSaFweOecP4ZY9Lx02huAH9xVBjGI/1sPlsIU9DABbUmj6I4Li
9hQnYoOIbFh1rAoMl69Qf3iN8CxvXt3T2OeDZPn/HbBxJpKcq1I8Qqu5G0u45VyXZBYNqJ7X2Ydl
EiFxxdmEj2+GG/vam375MyA9Ln+f1VAp5wUiw2QVsjzvg6hkEfXb1jHp2Dn8pnjqxSTR58xVwtrR
qUXctv+/ggKzotf18zTzVIvPJMyetAnOpylWiCOpHvYbz3PKTd9dwwqF6hFH8ICveAxz8elGrN49
l7gfqSTZEGZYTPW+Mcr59wNv3j21sOhmMwA49AblIEIu3HR6ClnIuMnxpdaMVOOCWP4zsRHbtHr7
sNl1jjFX4C0mihSsGcNwxJZB6ZJKKLwZH3MrUZngFdwWTcEP6NUZKYfoXdDkT/n+89DSvRWP+pA/
YGlkEzQnXvlVN7YsY9kCb8ZMJm1SgGx0mhW5QkDxFGRh5bcG+JKQMvDvGQLxEhkPX3Y1T9Jy0zT9
/l+0+kWiFSaus77tO/5cO6x53rQCZgg3ItuyBTHekOQFnilc+MiNjpqACD7eyt3EDfwVgC1Dbglq
SLMcm0J/tXayk4g0pTuGUxH2mEpevnd2HG0ht/vsOV1hFERVM71LRZGcSAxizwUw/xdRhJ5q/Ef0
auzsBuSBmmZ3zp7N7rPh67YblVP6IKQQnIb9CGo1y+Rwt5KgYdXf52s3Sx76C/GZFGCGDZNJDDMt
wY+lPHJRJ5E9cLudBdIL9hEMfXE9p4NU2UdJgqr88ZwGphOKI7awQt2kDcfsgdbgspd6DKIe+gBG
PFLZkwB2syWkid9WcVIrNcFMFi8npCi4rfEZ1UdgBDMIIrSNQ4C9KVNRYXWVrp93oIZjLKznZekO
ofOqzSxi8h2KBeztImTupvOzX74A8bS5ixZrSt/u1oRcIHsfnQSj8gT/BulC/KqlTfeQ0R+ZecTl
4eny/JHwKEqTQFUg4GkTae+YQfb5e4ATwmJ3D+RHi+civhpdiA5iSAamyMnKML1Gkd6pgIxH/lY/
yhp9iamCPzgfZ3y5yuiiWxglfZJc5bQOyUdXyuDRVVGdaAHOoUbev6+8ic8JGbbSmN0q9rRJiy2t
KpZ6X2Vt3pBgNiGSa5+UA/Scc1sgAQ9a7F17x5lht0kFMF/NdGY5bdIxPtJGS3t8O/k+3sz2c2v4
OhKsco0uRVzRD7qloJj5n71S+aOnUglVVeTKE8Lb6RhK9Ckkk39w8lGJ9X/JcDQNRak9cZe9MwE/
IE0Mq+I8ONBNkcD+6wjQtA0GxaUnBXDSpt10BFrYnS/Dm1iTaTF1Wv6kMe7sGincBEgArkKct0gM
3zDcGq4oQ1JQqqF8aB7g7aMMAUz0jbBAJ06dsRkDWsjpmbSa2nhbG/X0H4L1Nml3noe7bjBC27Mv
VEhF2ePpT2FHxg8OTFRHjWVA/raVyrJZ6saIKNRi9lOeO6uAG8C/gTrDuWtQM8MwYdCrs1D2XBvN
tL2Q1PeE+PAvaQZuDl7Xg6SsowjL0B0zYTqqN3oFfRmIVXIMoZ0LZr6w/xVkFMuaykW+sd9WA1d7
DCD96d0A3EoE8EN5oHhRm0wNOyEKVm97t8r0y3qabXfDzBL0jLmPakPNJxlvzOBYxxC2CTmWRe70
ppaot8TtmvtjmFTpw5WuTisSQfelTP2SbcHXmJUmQQoqPIDTp19AuqcNTOdtvP2bSiPMTTkvFvHy
APSXhty6VMvwFYZ0ALJPtjJxx7+Qr3sCv8EQ5/qZK8gIEREX+xYMNtxGHYWQPwFhfTaoqG7MELRl
h5jOYuJ5lBsJCrVBzYgN08JfvvRto8oWKzPRQHTbL9dolG6zw+3aeHyeOTYtYaK9iN/QxZI0G/zQ
WgQLr83YLid8HZY2VbGc/UuLQRLY9/TnXhx/AljgDvSVb5tYQVtNH6Tks2IYgeog3G1yln3MH6gu
o3LuObs1M5scLsqRwngsw8+UUTksuAkFx6RuvCM3wpf33abYWAiCfmP49r8DV4DQqjYnT+4IEHxq
ym7bS7TfifemYCKme8i7L/UKv+6ZlVdQoMcjkE//zvj5DbCQtpx9zE9pnFbAcVVlpDRnxE9VifS5
mLK4LdiPrN5XtmrP9VYrjL4edPSWzoosUBmFii8Ead3GZM/mL6f+n/JpvCLl/R1u28BDSHWf7V82
RoTAxCqNUS2rTUBwKH12rlCrJbHuZhh3I/UogE4HJqkuj0ApWa2OsQ0AZGzP05EuR3aJ2uu+N5ZL
huXPrEslmm5XPBLMIz5BBNy/ZYrlxglc7iR4P/z2g0Z6wANT1+bcCyU8gaTGsAakWap0Gf2WGv9q
ob6gZp6cpIOk9Ng0x7OT0ecM/AWI34lps4G3rj7d+r4ONolwlkMeg/qOlnx4B7B0d3Ji2M/fNBmZ
F2csZ3FJyArfFm2oj7aH5RoF9lCe8Z+MgOvna/c0FOtUnJHbkZhmHqk9zSXSbW+fE8Do7NjrBvyM
k4BkjpWz85BPxZLDMFkaYVzykTpbGkCJ/her3PMkRl/oD7667GZXBLB6BpBacsWaf7JoRIB0G894
h+A9Qw1iE1k97qy+2rbEpNOPuo2sjr4e/zCRCCUv4cF/KS91M08F5r52FvYVRTb1O5r/3A5TQUdy
Ctcoq1AIIEubcbef1QOr7ngqr43DdrVozX/vlPSqNB5CIW0VlZ6x5JSwRqAGiyc3PB+6uQl35r1/
s5H2eD1oG2iFq1OcCLr2+Yu4Fx/BpjdcE39VvGHMN9mSpKc1jF7Q9YGiDK/W8i8I7y60NcmtjoLe
ZeDJDW21Uez6M1lWuZGk+RbYFkYvaPqRDZBzcRIWd3BS/WXqFqX8n17YFHPgqovxGwevRSY/DBhr
g862HIgWs7mqOfb69zfKyhofim3wOWrk9bmNZR4KLTLsZhjlTX/zpKy6JJ3YG3wOWu6sAxCwFOr/
roPybP498COJBkD00nUwIf5FECt384FAhPkpQXyxhgJnOTjiwnApY91zNav45RiN2zB7vLcOqU09
eJUJezfh4lywzR7S6phWWqGEkg956zIq10bPVSYyrz4qBZA5CSCVmwgE/1pIYdvNcPB/3Wx+puaq
+7BJ8vicL2afSGI1EVvp/wC60sFfsB16Zoz1NcpTlyGW1ApXtv0Yt6964u8BEn7xrXRvdoSGpKtB
6kI24Uj/pE7G6kZiDzyRsWy6eOVTAqEet22C69caCplIad3kY7RxCEJHwk5elSIOp1PcALrK00EG
D2dCDdD4cQ1Aw2tGrVg4B6fnLGdJVwdiV9xeQtoA+2oeMbyVuMEZpIPSOcDrTJIOkgY4efAN21S3
6wljkI/r5/ogjvIwcWhAMP+dqj8+5YDXDy5CXmWePd4RfXqZpACUOgwqQOKYxYE3dN32f5zUowDX
vJl9PFX18ib+4GHA6hms4gFulwog5XvZXkZy1JAs63TkMFnZqgyIn5u3GUjavYKO75FWDQjRJSQz
5YIPdtSY7GdORjfamNE8N08klKVcm3J9gR2b8KhE6wrsADm3tnrjHwybnJE0Km0FzGDD2dp5trFN
ssO9dKvCMsDnDjU7KeQWioQbxfQSpHQtDZaK1He/zMeDExy5u4zJJWVZm1JFyGmsm8elTBobjTyG
heBvibougyAV4lnVcUeJd9PMR8lSoKtEQXW+M9DEFCHVBnOv9wGvUrshZUJ02dl51gpcASoNE0kw
hXz9U5PpUroNFy8z8mmX5xHmTw/SzviaUMv92vnhV7k9dktUvQCL5pNuPo9R9xAKFfs8yhnYDSPR
GJOOQsKlVu5xpPgts11npKX5DgoMyVQgyJSjr+eHdhQxtBpG3jVaGvtFzKMCAqcK1m1bfpKA7NQN
CoMNd03a30cfWh5OF2cwzpQOCXecfFmUKV/xqy8ZXt98IOYb8p46YCc0+TMqCTrBASWCh4JeFpRo
XDZdAlgho4Zkq9yXbPjy16OPb22MyodairtfYNHHLYAtVIYp9QgsgLApiyfl9ernNKEMt7e2PXg1
gnfq3FaiEVVFS/81VXSyg1bvbxegY4IUhtOkJwCVVsYiIo0epomj3Mm/9mpLUoHOedtGUJFtrCdv
i7D1R1M4MnhRGi4i8VP55/xFFNn/IiyyU+HbSUuYvDwUWQ9+uHlVkqNNm024ahXYPybY1o7itZZi
+gmsEu6Y6N2pXTIibG4YXPL647tv2p0gOqNG70MVFYFn7UaZUITJcd1fFBz+6TK0eW5NaMzp0ylR
N0ElHtXXgbwmHbYPCDlydkSA5e8pGe67eh0VTHeARDo6meLOLqgDAhNv9Jjz9hYMp7+bzsgkwOxG
BhUEGzOOkJHPQpBtqoTeUBIn7/jr3/OuPPvmhOlPTv52iOWuTq1IMxq0b+NwreGkG5XejNNi4vvW
7IZF2Hg5niAW/sJrUyV9YKZG5JcVGIXnhYnvOjPDi2S2jd6ch/wS0Kl6QnskaP7OYr9ux0bu1neZ
ax9F55B0UuX0q90qAPvxo9XGRUS/ZMBpJd/xzA3pu4Ud+UK57/KRkiCT0VxwcYwZw84qcDC5E+hN
TP2a45Io40HSO8/DJBfLQ2JHwSoSjWiyOHKmjEMmQdA/9dXT5S2nH454e3A9kgPPd7HObjsFEVlX
iCc8zs72RPzJ+se6cypL2TXDrYJJaeYkog87N960Yl2aUXvWMfK7aKEomouXV/rduAZo8IENnKOl
zRGHvU2WGXOiMNnnnsLykd08q4sBg5sCfeg4F8RBfyshXDrp/bCCx+P/Ajhyqi6xG5ijJTiZX9GB
rMOMav36yRGPkw9dUBad6fzWkxVHDaAg5BTdLpl4i4OqW7+Ve4vK5fPpmQxZ+osjyhH2UMcFujTi
QqTdYZLnUqbUVtyI2SF+kOVDLDk3TNdXYMxmDudvu1wPhrMtf+jQhlRvQmeTaTPYLjZbNv5uNkfA
WJRoklah/BxFmT1cf+L351GvHYDHW3Jl9k2g/ZLgQpDHOWhUmUvw5wjrnNQxw07cdiEmQwaMz7Kj
fhJyxDNUGeApAhupSkhD62lSe45FVvKRCJPfRXznksLNzIHEP9Aeoijz2fOHLXal9PwC7a5fiNMK
3MqRqFMWu991wnk3tF3j4+7c8iyJnhX5BlY9fIRR14bPrMSAPACMkxENdDH8+J/fs6PEIPtuu2ex
i39ENGwlIgd3MPLFk3WPlxCJl1W0P17I7OmRWev0ItrnWxdj2DuwcqEefwXOoiAWze+p+xyJwMQ3
m8HMV9Hlg+JJEpUW+44Boboftfh+sS7nxAOougBElM76jbsY+VzPczoEueav2HqiP6NJRwsMPl8M
bUGwls4DvCvQ+r6+34Nfu3XOrymHFkLljOkHWt3Vps7jrNs/m+WO6MGDFkOdO4AXe8LCcbopBl24
LeYy0LIjyjYLjpsJfOmU0jdCFD0SJlbm0LCm0Xlc59mPqliaQ7sfp2PcWaXuQcD1Id4mDWQBxTNE
RFd5CpYE6UgvDLAxykzz+UE67O/RwHBhmJsBh2Pl+RKzplVnu3Iv6tQkTM8GguRhi3oVCd+lL0H8
N4CTrGGogeeu20mlPfPa5fRiZWquPne1ckMRYC2Ze40vhmicKCYibPGmjCMg6EkQDNJqWjig30/s
5nQ1ReNwlpW62QcKYQHiwtwIr7vP7jA/QzLT0i+mH/5rFyjBaggrOoAQtKNAdsk1yHdFKw5U6yQG
CDi/rEviVOtbX6ActF4TCaJZIkG2E5uU9VGk3nKhH6QboIMfUKqPHxyqzSKDbG8rg6QiiCj9pmM4
ss8bEDJC+tFHWbz5sk4Rh6GJdb0q6KLFXKdTrEeDnzRHHRm4D2YrAkWSwsYAX8lz4MpDZ+NslZiu
V2XP7WMaHwqYBEaKuryQnZnVTXz5ROY3Mg1rASItat7x0xHdzI9+rtz9vByZQC47qn5PXfeJh1mo
3k/sAkWgpYpkJesOspMZjXBmuvyUdwrQTyzrOtwNkD45a/u/IUakxtBkzTMM/SgKwQ/Oep5/7W7s
k9bH5g7zUM58UDmeu5yMELFW8IamkbJQ6qtBuy2wZzYrELLaOIiK5lc695UwnEachvKjljc0unLf
NOAHoYCejnrUMH65qOYdmeksTyf5k1P6ZqM95ouQc6Yb11Rcoylg12tLt3p0KiMD9ZIPR5vuWPoQ
RRBkdWRb8Kc6tij/BD6ZGsFTr5vyJ9FZTfOD+0C8FQBkpOlYCjn3u+I6CSDXcP+pAhjRM4LK18Ai
khYxAKCanEQ0V0XERDjel5rye35LRfMKfMvXp7lf3k/einMndajcjEEeq77e4N7Yvxg+nygTcN+m
6dVXGtOtzawEx2dLHsBJyx9wXnlj/QeuUkzbkyxm4fgtjQYlPB5m0p3eSrUmjtKn/+Ut38fskfdK
q65OHIeiJN3sBvkwOkfcf1ql/izqUVAAVRrLPXKvzl+xNxDnFj6lcigiBbNScEapeKTIoRWfmINE
e/KY6KeacUmxC8VNqoHttv4Ul68MfJnfmT9FhNNqqNjjgbYfkLfTeix7tzT+KHCUJQpxFdQfXITB
9F2y/GqbYRT3QxF+IqpaTB/+U5vzgegdTi63CJ3/vGs7fOrgRtxW9cm4RDaWK26UYQGPt0VJ7+OL
9+KSC+PNTRa+7jl/uY3eISv7Z+Rt9koH9D6RmQUQk/2MowUpT+mVdoYjIQ25+3abnB52SzyLHvLp
riqRPI+9hbil4gEl8xzouv9AgT6fxEfBfgROkfsWqNoDU3sBIK3FOdQdFWJ7GN4k9nkv4C84Ytru
oDmi9CIV/I6jpzVX50+F9Ll1IMjRAUGDMFyswuEFUaIHxkItVdBsB7oDc4S6bW2M87zV4PxCq21H
1GY/S4D7VqN4zc7lA/EWZIdmLz7W9WRHzZSEcToySwyr5NGBNu7pEOhdbqZX7lZAbf9rJwVAXuQ2
boJeSad12KJSwahnT83o193/TwHJOtK6sk9E6jnRCTzfvi/vbGbs+rpSy0buCUTqdYZC6oQpZZ+Q
3BZEiyrLbfcrA5fE/SCeHepHaLqBBYThrQsgSri6oT31YOsoWi6oC3B3+TJaIW+PzaI37m8W3GTs
1tEntl+l9RjrjNTa+026nS4SujjXRQJoondnxVHk6TeT0hlfbPgmFfSKcjEsZFxppPamV/BMj16s
J63i3O3ugmz4ubqD3t/Vov+yn8Fjc7FduCPC8ZSiGD/U0IrtKZRZ8+c2wN+XaSGjWT5XBw5l5uTk
2HJFsjfBxx03NKsXfxQkWw4p3cAWw3bESVoQu4H6FFfbbIO3rr8C/WZKvWZkQPLs1S1Nz/WERmQx
tkqXpF2QhXsaccpn/9g9VPqHouzOnzm+UtKjzuRAK4U87qKeQ3mofjCLhg1N0tya0OziEsqy0me2
3gbymVjnaUv0MeKrL45m7XRD2A3mLPohCvGVgzl9dilnuQj/wBYmhk8XvBEfi+Qzt02pQuwDWIeo
h3v6LNaursjLsJQf7zlaHm/AmiAO5q6sS845eu/Sn7gevqm3X7nrnAtYCX1bSxWiI7kfunxHBTWX
02Nyp5lIQfXQrxwSvrmGKi/4It6nuOf844HB1knQ5BhtEgldb1q9Zo1ygwaJJ96xsxi6apUX/NNu
TfBaTbq1t8E9PMUNXE2Xl9kqFuQBdaLa4ZXCTL278eDrmeYiM5FI8467UKDFZXtcpqQg41azXG6H
fV7f4QjgxlgKNXYaBIfPCEytdmAmSAfKTfAWXQ6RagHK3FxwLTM/wQmHfed2cl/BL3f9m741E8+a
DQjF2QDbe+lKrKATJPGHDbNYwGwG/VJ2fb3b+ZOhMVyIjmPKkIU8KKrE4xMMPXJ0GOV47xChz913
1iUHuK46Plv5PVJUbF7nXxTgXl2uVE8vbjR+itFaMZuNV4taNG5P6fTPGsnQrntSYNOon9NL2taj
HMV5dhIZvVUv2iXY+9vWnhqu/zwBIJemeTNvl0sbzym+/Dmoh7mgSpPVnMK41TiQFgXlwmlm+Ec5
UGFmFVDWt1gwufK4HBcKkE4EQTC2eRzPWi8Xpfoivmb4orf3sFeQGRu0eZu6YHh+JVtZFQhLuWFh
80STANZ90+qL7HLiOD4v+PtkovR5AtcVehp+ADw38nVPQAYfFwklBoakVG82TU+pLknfHrWToBJY
Uk/hkG/jJcVSIlb9YIB9alUcTsBAZAe4So/t/XnLAhrV6S0ZZKbyEjob9fCYpnwMxRuFaoZnkPQM
fT6vquPLbKjmN4SczE4DpcwrB19SPg1FCZOTKDd51wrLS5S3qOUGdmiLmSV5FBYDQ91lgVFOr/zf
zuLHQITU2Y5lYyPVqrFc/xlPS0k/JT70USvnLB0RZcY5AGO+DUSdjCoDcEw1Lo1tpiVDB9RUwNkq
u0P2z59+KUAh4Q5OGIu3SOFcnqKB+mm5JmMBw22rRnPkWZg+DedqMxpluO6YXF8ZaSxEugaU+nJG
t2uOb+mpdyXLoI8neQy3eicX1QQheCpLolvs5G08bvn2ikknCniSNROEXI4+khMogQ6U2kEokz07
xoUgsh70nXlNrTCz/IhDfZn3wOPeQFSAV+SuQqDwYVRPR30wDmSHEjvhweJTbh4nFw2A77iQbGEq
0y2GFRFYhTnlAQR80AwbejGXHpjI2L+c1ppJXHPb8pP42K9hfml9JQICRhjYPLm0dxZWCW1IgV4a
k9Mak8jVCn3i7iPflIQYBiAraDCU7uh4tKq33jfkoGl94qvEmlEqgGxXPBZ2dZBvqPaQcAkh3wnv
Mua0+5rDfvNOrUru9Yjb2r8xhzm3U5retBA5we8qF3dgAeSNdFAoKIOVNQGAL7JzymPywvKfSq7L
k8vSms8jbxrxOf7wuAW86ZMfMG3Lluej37gyg7UmQMN+abZDqK4RUXo6Z7hnA4SiwdVzJpqXhmR0
SrZc1ttTBDxHQyKQV9cTK6CC59BWsHhuEXS7Ct3pIVAUBA/R8RmLRrvihlTzGoJg9Xh0SRSkxQ6u
dRXujWHN8HV5urJtGG4NehUFQsl8uPqCj6yzsU9/MfUiTx/hwdnf9beyuY4jEJGy63EuOGM+Eak4
9UPT4iAOXa9e8iXeqa3eJJ3eMLxohwWb13w2hXXUPz80pHC0l6vuyaud1o3YkwRZHNhbf+qQIqRH
mIp6xDzOC/paFpbjCjefkieWLzgexcliyDMEIL/9V4S7UOPMVfUk1UqUa31S5MC2S28ibajfvni2
o/gvgXXQS59Cy7qxZprfNu3qe+qQKeaQdlQKvHLuwFAvyM+96JlymLlGJtyM+Npc2sWzQ2YiiL1q
87lV9AZzD3OLHBQ9Sa8MEtLP89wHBgbLh8hpPTRprNYu6veg8a8H/BklI3d/vXR7pDEkiUltX85O
EQVtcLzidG4E/wyHc8uMMEr/RQKpGj6udcF/MduL3KJLputEAfuTPZQ3KbAWsts4i07W2BU9AkSi
Wzl9PVE9HepvD6eKJt58CJkDhSAi4EsxDxkXlb6ZrldJQZZv+J4AMEFgw++kohtmcy8lh0BHBMNt
J6f+hXnTljmiu0RJa0PzhT/FAvWwPEnSboVhskthaMSyokDcIz0TSf8omnLG2z3xJ79r7IL+uvrB
g0mmkC81rDRdg3+bTaHN8M3Hz+/ZtFPJK5EB9srYOJE8MKRIg+oUtaN/fs8bONNCF6dPzN5N/jpt
fakIR+qmZL7Q4vSQN8GO5yRJa/oDt+FAmGxCQwPjlfg1VMq4GUbz7wV/crvRZCw2B0xZrfsbqMra
Cj2G8eU7gSEHS/ECkXMcMKXeZ2QlG/o5bvWlKzr8m0D/BpFOYFBlaNLmIk/UuO8olMK9s2HvRqAq
TfFrJdbnyYgAgvGn9MTiwcoDcZ4WtS/LuMoqh1CuO+YUzuHUSnIhpHoTom9LNkY2xFg2QsGbpZ++
++0Z9f654PgKpSOo9OE8qJX5qEaRBXcPyOqT37H1lixhKTxc8DoxYWFxcHOFjKdj34wL++e1/pJE
d1OvRhGaWlH59HzapW9vxWmCm+MZOLL7y+utumNWzBGp4Wejaivqe66AJulaKAxscstlFJTcze7T
DYXMKrrVH00A3nTRD5iGPHIfqNTSPYAYAES0tXp/txrlkAOtKQ4LnMy+c9WcSHCJpfVx7sz6JHTQ
RTrXeDcy7gTM8YmTgAmAHg07FoxGRti9NbD+CJi0StM5m7FgK3T9TGtxxDauXLrlTEuWRfd/0Zj3
RajSDLat8nlxT4bbflCEqpYslXHh9HIvahynr1pk2yB++sABB+IKj8xiT2lzdioFyGoW9Qe0QFPS
YCkATmUgFiA20ZcKVaGjSKVj3UBdQWqjGufdRmoSnr22Ums06Y/UcXdE5/3jsnvjyjbFjlTvm6vQ
I3CxBy5oo02htk8Y22nPzr6I72BLkd6yTq1z9RacdedcHzB1j1I+uNruxyRF7UUFCKHSYyhyGvEG
0Q0TqWSZvY8nRjimDv3zSanNj4DQ8U7TF+GQ2gyaeZst0uBWlZRvRKjndF8SFwbwni2mF8iJlTep
w3ncgi3FW/mh7poBwawslyP2/vrpYpq4kK5SL9N+l372sRjMS1tqCb2e9+Gr+xWpGbmvmXZwuknm
IAfH7eVCIebx/iOYZp1RoHrhKCUDzQq6tmhXsXhBbPfe5xzvPc3F/QYDeYbe3x3UIfChbtlp8QQ+
GA8z/+7DKofJf3uRYkDjyITv1z9wP+UCS4HJpmq2ygvY4twW+M+Qu164CtUzzyAiDwX00l9FJTyV
DH29jDAeIRuxEwqAzGK7HuR+8Fjx7A3G4fq8JirdOYpKUOKDgImdbJHi2WbmkIQ2STlv30gbr1N2
okPJIQ7mUid/2w5watppBB4AXCR8d3SifHokoSuPhOomdzdaX9L3BHSsWBqjzaKJu2tewpNU6JPO
XjBre3hQIkdCWbDggo60tL+UFAqNCAWEakvKu1cQiOfRhYbMxezOq0g7uei92z/KFoPpQsRohXPS
bWICH+F/qN+WtAjpo/CeYjZ/ClRSpkpk5olwClpxBGDZdS4Y4y+gFsO4SBM5FvDfLaPwLTsRdBvZ
WJbjioQPrB2nMevpc8JBuGYtGc9gNaG7YhVCd5Qat848SB8SskJNh/mmqoNLqeSbt1zvGmPTu/xM
+NDdjVG9+X/SrAHRNSgmi9Y/2/421mG2Nf4UxKU0jGiGKGTsY4yUyMlnLpRm31UgrOlxRZJh899r
pcQm0wwwGi3NZX8fcjJPZL0Bz6FycgkKGUvxrL/My5HiomtGvEpQwVA4Qp5h3y2UiX9yZSW/uMTG
rFYOKeKcKW/Lf5Ycns7nV1CWa+dXyytC44G1nMd+SkWVZAQstD/UCWlXy3FBVfBjeBTvJhMJtLU5
r5+sXvOAgaoOXXp8SSoBh3/4t8OLWQ7hrKmbRvnxV5DJh60nWnQ+yGICYsu+QQMP4kNogJMRec+1
sMpBavxiLvitGXWWKgG4NzOnGHKbMKNGKQ+Yr0di33hES6kWnGJP/mt84gROG8uATfBBrOuwVOK3
geHpQocVuaG9K0/JB/4BNMcdpMfaC4D4DtBOqtDQ/ILIOL4ZWTh/qlT0NxvsnKRJbx9YiP2krvqU
ofsX1keyW8Tt/r707kCMIqZ1DA8uU9xq6eqFwgVnXQ4SPl0vnSc0wusDkQErPW1skfxkSj0W9u8u
i1L9CwKg1jUwUfOc+VUOs1OM77CiqRZhcccn8x38Sp1lYPzPDs6ALfCsHNr7LaQbQJga9Z4dol0v
i4kpF88n27CCRhQnHbOwCAqyIuoD4KG9R3tRNVRYWYpJTh/DHlX5jBo3n6l5n3UcVHv8gqv93Qbl
DyITgMpKbyGy5O8czJeO2CHyK7q5Mq2/AQimbhxSRZW46uqkjb0ixKMZRa47b/bfNuMFB8wkX5cl
k24bw9o9WO3kUcab+pqRYZDfyONkttEy/oFqs4sVI2JVJoZo9TWirfLxEvPKolxFvv7/9CoanTDS
DENG57hc+m2YyXKTqAnnSzwihsdrUoRMZ7mwV5nY5g8V9NwW3FuA2ykyod8tn6gfb7A0ds+3j+jx
/y7XRhyyu+4fKj5Ze6T7/KSJUx9l6E8y/sgSTnOITsS6pztUVZPQtw9Rf2Xqh2TiCa9Lgq9c+Ujq
XoG+Lp4txk/oi305RnuqHN7NzBA8ce/uKzI88ClraWU1qAyL5+Qw9zGIKyMD20UtlS3UGNTsK6FX
267I1nI6/xGpFDmpZzvP5EjbcuJ0EezEqi8mjtR75ztsnes5XnI6ubU0sEAhJSvrA+EQp7nTlHG9
zjB3U0CKyljdVibcbSdcHigMCCoPkwOrtCukAIpoms/6bYfLhY7zCdEWlifuOM8OdgAJ6D2WScVn
5Eql4C9RdKi8ZLCjW0IXsgacqzwO/kAmA5JI4PIXuRNp61Bm6rDEGmTOWw+NDdUkshBrQoRQWqhF
ujoNYpJUQZ/siAelwPEt08iEv/3Ys7skJijwSQ1oK2xVgO5xBebQJpCL5lx90jN+TRbrQFATf0YG
tueY0AOO8OKJiIvbHAx4etLVpjjeYIt/ragU4dZfQZJUKX9+AIFSbVOdZJg/GR+8amhGY9HoLoLA
icq/Vn0/KB26ndKf2jEnxF+DJurs01BA13AwOYrYONl8IgoHT4KuXMP82R16PfIakk8jaO8lo7Pl
DJ/i0f2eArwuJYno7SYmPFVmvRrvUPSgvXBW4mwPfWr0tbjvPmPmFAbqS7Q20iQVdHPX7aG8flOW
XxyZuUrNqS3FbCb9sUvUt1/FYyH5TVKpK6Un8TBehFRG3kZxF2Q36lRyyemJtON455ry0G6PT4S0
68RjotDRwH/52De6WH3LsQcEVgKo2LukTg6MOl/rOFkRsAIVcMmMiKexXZdFzLmwBhPMK+LiEaa+
QV/RLZuGVH6sEEuP2l6IWzSaY/hSj2uJUB5PGTUuMV2A3ahjGHR6mgUoXsr3ReWIQesSbwJzb2nw
I59d2q+V5Tlg5CoqVpLgyxrOnijcZ3pRGrLehSkQKCemvKKWxQaJxzYNs7lLc/OcgLhbxhTNN4Sx
Ac/XHZffnImJLGOJ/ljDsH2EqI8WDT5V46EJD1WkNsbcdSSTQ+BXtTva4zsc/oJvI/OmtvtImX/5
6HMazvwZ0kl3Y6CNpN8APeBf6NUNvy7Vls2OdMb9UnjD9qlC7ZsMaWPMXtondcaljYTUNd7tUSsY
MVKK0UZMwS+QRZ1vUSnwLqtRB7zUh5wLWnLV/uMNup+Q6S71bCATTHk+tbQnSTvckKJYy9UzL4tD
gWDdQUG5QMwo2D0AyX6f5nfz7E+xhKfIOKOsuNKMhVqdBV7YPYVrT62Xmvpdq+gSniKQ1n+hiCkr
SMStDg/Pwv3BR+zDMqcecv88ml9tjSx7gq9Q7tEgho4LOsUu+06F89CaqsWoe2oKNn0HgcZ28PPd
vFohp9qsSgwqqkb8GVB39XVLw6LNmBjaFK87f+bWTVrsl5F6xeXpcD4wYhhwEsiFrrvchXL1pkSs
tFe8jzs3O8A0iy2lMq5fj1Dpz0+eWlE0BfHKQzYLY3wdVosQU2kcDRbHe5TeIVMdqm0yE03wPzp1
Bm2UgfZb5nR3JdPv3H1HIV6cSIQsk4S9Rd/9tZ5CnZqDy74/Ml8s8ZQIKDE1XqspRF1YXYhh7lma
fVUCpmxjJfiYOqmQSUJStyPFsfc5NwuTD/K4S/vKTo73Jw3gLFTo5Rcv4OCcaMKqoAB/0ShU7mgn
QE9d6ArTxhvlJEz67iumBdcvaSjU9wSKHHJnvfzifEx4kLMeCzpGD+te437TKs4K4kCYebAwvM1p
i/K1rc9c7n008w+9BgHSQGfR+QO3EL0qfE3CVhDU2Zqek9iOauIHbaLsPf0zQnp3VThZaI54N4Qs
JzVD1vT4cdJDQW3mZuUUM5k6zt3KZ2ydBJ9lyMUCt8bQtrXo6diFN+BtBkG/fP5ASrYNbQ06gLoc
iXfXeFas6BxgrxB4Q5FBkMyVu9WrCq66TTrS/+dB3o2I/H0v7ciNuHqHJAQ4vn+0keInR/4CMiiz
2r2k4EJnfz7vx1B+fVyjo2uJ+U5JRhYuDgnDm8qX63kSvDo/ngC4Q06wWYgfJKsqRQYVK8JNWzr+
yQ2BupM7D7AJnupaHisjd7QtTy0w9VDbYJM65cTZfYT/xx3lVT+pBEzLjWbj0tsUhzesRVXmOPNl
P72bJ/T0KKMEVkUVbZqTIxI0dRRcWsO7+cijq+ygbR3N3pN665omwsic8b6G0rY/yYtQxf4g3S8Z
JAzH5WRzjxlPWdXg37OIrEeNic0oMcrdTnSHnmz64BvwRP99p3sOSqj28e9X2pQZKxsVc0f1MdQi
3cNnAAkRy6AuT9xqjIrVHEF3bmS2p7GyTS1Iv9/wI9GcKkiZxydR6v2Mhwea+wc1RcwB/b+t8UhD
e+CQ5ohLCKak8KM93vY7PHeIETqFS8iSl+Slraliw/5fnGYhHWcshBA5Y5+Orv89GiyGOBhNDQ7P
00YOSpBezUbgcnitqjWnkTLKVZpYbxo+7EONyenEFloPKcr2R/ewvwnzkkgFBvceFYXZ/TyqX07g
0m40aniaxSAlOvUgpYZRw9Tcu0NBxSuO0L62ovMwvtvp3yXbt/uLS+v09f25hmdmF/L9uq+5/5AJ
dIolBlKzqBBa5brNKBiPDnSrI9AyOSXI02HrXWcQI5N5lWjsv/+gFsNnw6WBsHRteBMhgdkG41bo
L3a/BlxpDTs95lbTSZrPiRp+3A3y7Y1EJSjoNnn7fvBih5zX+7Pqctouit4R+lREl/pKpwmhFRX5
sZ661AQtgSBGg/7g67YfP4+X2bzFM3ZIYBF5APco0y49fA9UKWfaQ7ZODUUQwuTEowB7Km9ivTah
Q73YuLMjux+FmWaq5vERNqQvke8mj2hU/H3S3Fg47zYqAfKpPP2lma78OjzVk4NMesXoe0qklPR+
x3XzQFPLjPod0mYqZb7kgNhclaa5Ni4df2GxQ3Mi+USkKfN+Vpj31VH/Mcd6m6CtcZpTFuH48AvJ
jh40TyeJkdaSpwGUYrM6MYoVIMZPmjr8gcjzrWvZXqfO0btHJ405CmhoU4T9UptI3SrUe+6BsNK0
wHMoTyYOYp4/AA/W7kgfUktt45DkSnEF2gBkvAo4Rtqd691xdKukbB8LCqx/Hi5glO/DqqyGYLKG
1eiolhI1niC1+iTyb9UVt9nnj9DT4aOGsidjQL4NibYI57BniYiNvXjqnej3U+ojp1ISHvaIl3/z
47bvHaC7n20Df4htFFJzTWMdYRtHOXT1TeMPCaRsyBBIQE3/rjrYtYnv+guFOq99K0T39L5DXr1g
l+kr7TvvtioyUad9I+XYaVik3Pb58MVfH5eatz7NyyoGyNusd/bnoq7epe6nQPaovoaDtXI2Bq7E
wAQU/jmyfHbszCANIxRYmVARQ0ADqcsGWlx8iZhT/OkE7bHP5xB/X7FM91X2iNICSp1/11cqoCmg
Z6eI/t9ljNelzE3VWCnI1+5GgeBR2YGSAJ0Y+82RPjAUDvP8y2wx/HkLpbwEUC0fuZ65Qz9pUxSk
2sjRQSzuO9+0SMKwtC0N18mxxhrgr4v/14qvc871FGiR+FmWRSjN9wRBuPxbqAjeLlOSu46QEVAV
PExlh7zzUN/3sZE9ZH3kBVAwoxYVkoA54hoaQqugn7kHm51CPB4C+Kqb/YFpCPhI/r/rcZhsjmvu
NbFq+f3miMCyq07rGVUZDiuk1d6M9ZFo9J+bvtiXzV9HNxrqAPoS/1i9v6h9bMexqg+bI3Xam0FQ
nBMvOq3NAq29yo8F2COcyH+12QmeyrkOg792bKBqsR4eIZKrJc/AyTVxVe3sakPEQQkJo5byszbv
V7szJ8mc4zuki8sGEzgzTpOojeAnJWX3VTA1WgE9GwH9epRqAwo1P/75MC71gPppQL1DN1s3LFks
no3qHW0e9/iTzUomGadUdaCpG/+Wif2MjcBlJtURcYdnUQb0Xgv41ruYFEjey0/gObAS3gpuJU48
9dwgPYOPnO3oNH49sMgFkRgGWq0XtRsw6WtD+WzVesLjIZEudhQUWueBAfJS1BkkRXolac+josU3
lt8GNlAf4KskYbLeWvj6al3jc9hHfbEt+rTzWxUsAzOadpo3GtE0ZkgLRQAH8pkC51G8gx7KSD1s
N4zvM4rJikNF8+VOmxjT53aHYHcbOVY5G5ggXBfK4bkpPI2Qt+JpjxdkWw+gAUlKJha8Ebc5ZGpr
RYFRElUwVf9NEHLnqtnXD5YC95saIwVWgk9Ht2xIexm24OMoxRUafS7tXlJFOOcu/oF5WnY2IrEO
9eWM+fu5jq1c0D419xD/uymtxf8xmn2hJ8bFBn7JIA5hF2JHeQF3yGCNQUMOBbFOx8wlfbxU2+Yf
DuU5JGKxPFKX6Iws0r/1gbFyg6TWHRjbIkdN3YvH02uuLt/KaZd8emRdPxTid70UebdSrNMF7/KY
XlPN3peeSoEP1vzDpasyElULfL3buHj0O9czDwTHNtuCy9SCPj6Sfs+pGPqDEsk+T2nDXDfQGcLW
eJ3RtCY7kmL/w8uJP4pga2TiOyoaJ4LzEHrRmEZEzLNaw8s9D8dQvXW1VdpgfgkuH4Nn4FSihx+X
/FcU8XCWUwKkfzi20dMMbmK7l7Zh2o844v7I48E+MZo5yzSrtuF+UXGhcb+mIYIjcKv8fSUmgWuE
2uyxBQDDYeYNw3gqiuN/NN/R6IlrOANS9168dbSjUZ8giowZwolZ6PmmIj9kqLv3ladrFOhjkr3t
EFLAd2K4JCtOG/kaDZHRsWTEw2DuO1ORzbmMRQl1Yh+fRVVPoreZzJPICqmvneOZbBIkXiitBFlM
JS9aZWSLL0/eL8EVBFdzF8bH0yIO2LAmCTveZrYZkrR7AVq1B3GkeLPdEIVk88sLEAIjHfYU8TKO
luTnIEVLPxvFiGD1Ux8KAqSo8gFLQSKfDseT4AwV/QO4X/gQ4nVDOsx1Fy0+9EozbjxEMAiX9SXc
79MO1tgs+geMYQW61wKEw+UX7OeVtBNK325j4gkXCUpRMKWgbW1xHrr3/jzXxkURCcWRu8LZ0Pce
pmVzece9u5OTVilbi8C8MG6MQ23gxLCIQF3PmWOiCVDU9gDcLrbcHx/7l4CwmsWG+wOAIEZc9tp4
Ob7z2JdIdTDNZAkKLCAGq5GpMvOhW91nkQLGFUmvdcCsRnte9hbQ2BDc7cZ6YkmlmsQgf2m6Ns+0
i1W+EhjufJwsoJTtBu8wW4I9I9LvQ7Yc++I1Vp2MoeuGhsnY6B5LAS6TeFDt3sSxOvPP6DVcWVQE
/dszf+6doXfSDzWGkHIMsEgf5n0+2HqleBLEUMOJFfjOwB8Zrm2qS6mcgeEg0sygXzeevwEDoj4U
LNoe139/sIud4eyT/u9UFirtnWkzqrK804YDSTH+HQ2zNatrk215TuSi4pkzVe0YBeSmgoJh4ivF
0iYPLcHeInHXGaXJ0ec2faZxAs7XFwzyS/kgTsaa55pfpF38enD/APhy/E16zpyTC7WxY5Bgj1x2
07L4kUlFskHyTcwIopXersySl2JCp4aKe/HjKJFC/RLpyt4E3xBAG66hzlqwXoQZEgMU4F8e/E0T
DALUebjeacBiIGm09IfEas9D+9QYu4Vc56cqyjS/DHTfzL5TDwnDO8FHVlL/Tq2qOVFLiKsNMudD
o0sfkd4zYGZK4Hq364aGdJ6du62i9eSqnRZFV9Mg8Nnc5PsF05QRP3QuOAagLOMFqsrDfOBNckfc
It3kR/S7ATbh4/alDYKLJgZ8lB0zCXK1gEkXPwVdSzZOC6tdXfvBQt7j83mnEYjzW6t2+P/4Eou/
ppI4czQPovcpuJndXICMIOUTiWNjz0fiddgvC6cRIVeIis+30A4vFyr6CwdQ8LEl+MfKUGQSmLgm
oHrL7L5AR5eycNuwBoVGoS/mHj4hWVtHods6wCyADf/Q03HvLD210m/RNhW0msxa7eoDcQHatA3M
NErxlZkuLZWS8ljvvpMWfoK76Gywv2Dvsbsk/3VgMdVamsGChDjTsm/YQPq1ROEdJsA6W3Nsc++l
5dkvtRXgVDqUEGRVwkTsPo0Kdy65Er6/Il0iYXDPQl/zDO9yTrSIykrm9hqv8eJTUO47W8AjtuAG
q19A7coms8fLYZh/myZRYDcCLu++4pm73b/4LPLqeMoMqYGOtUf1amY/thL0TxjL5vfEXCaAUZpt
u78E1Gm4HjN5na3cgB1xp51bf71NENSGdyrg7WUr7EU9suZUv0K1QSR43/ZMAuogvPpMvzr8jhqL
sSjb7IXHYs/9df/DRNXwmtluBZdgW84+dJFN7q0MulfJ60TGhGLhX7ef8z3CIxp5IcA6+zQkN65E
gFK9SGhSkMKSWRyS4AZ2I68VP2ndHec2CJzCXldWw2Aej/oU9JH+TAiOyiRUz5yxo9tbO86Hpj4Q
vtcxbLplFv5GY9k1rWccMGIoXjbz8vFbGZQhsh5CAQSGWJ7nncwgSxcOZ1PBMkRrPtrooFyyrcKn
bSH5QyvkP6WFa/1EptA36bUkHKYAtMLZEkaJUR0guIvME7xrDw995llMe2J2KK57EpAoE8rFo7E1
947pOhj81GuTlV5QMkIMy9i7/alHiiDc8xoC7jHudvrQwSvnU4GWVmCSOq+TbstRgIHIjMsA58Ao
EqC/8ZzG66Gz+RNn0ECMUiMK7F6nbn+5cBOR1ck168cwYRz00aiDFAG+xjjguAnG7wBUhp2Me0ur
nRbvwau6+3s33LazxerBBw+jNhW/p/m/OU8YMfEkQSa/T+faSKjhtxcoK2bxXl+lidK8/YIwHI6Q
5fBWOBFBI1dun+bUg+DruXy5yUqEVmfgwt34aTCiCuDPZbzulCbKgkT8TNaAsYUfdKGr7bw7lq9q
rwjfPSJ7/wbewD+U3pAsE6+tOfqtty5hXS1QPWmWdslDIHY6qcCQr3GRcLcOC/VQvySYwA17ODe6
OTOhZfQjCIBGRx5rvNYMHST1jSajNYWpog/qso3mwPYTmRQA+N06sd6Ac3703nIVNF9xlQt6iUT1
MQXF4Hns28H8DLzDbyv19qikqGN/NVq9Zk8uNWywjNiYWXdOOQtn1jNHr5MRKYvyN2pN9/a8IxQO
Z638uqjXcWX72U7tpQhXk690QurJGZzp2WkGoXv/UgJI46J6NLBZhSxpsc4YdAYGtIRA2fVzBfF/
5hsY2B/2vZq9dbFl3QWmWzDHxqn71ENaRwTo4pPflOJCq4VLb5pBgC/3pmYny9lCrciKS0pV8IkE
iK8scS+ENf1+bME+3r8jMj7zQOamNHafHe7MjI3Ks/2jpLYemXrJUJk5+WhGIz/13iFOCMijzu5A
ZoaQasZOQ6gDLzc/P8DB2KxOx6Amr2yqBaNHFlw21AZfj/QhWFUFUIO1W5+i+YeLt31f0iLRrXKS
gpEh9kHWxdetRYLuCrreKM9zNoX2JTmkd7+UlJsyfF9CoEBCq+rwpnHHLyF2r0lV+d4szXHI2ZEV
S8rT0/exNmKpzkYbrjZ+N9swbhw1xCqov9LNCe4oiIeVaRWQ2U4mPZm7k65Wv37fNtjHzvaV4nfE
odiq8bLpQ97s0SxAazQGyEd5LntPlGrGPc8CshvmENoTReFk8VJaC4hlkC8wRPqv6Dm+f0qXYhhO
kR8ikZKkHeTYbHF0sFboOVyYWYUjzbq5N664Th9/RRqGvlrk43Qi9dJAJcw3NmNxc2BRw2lX+RVH
3Iit7MY7S3N0tOw6CoCFXk+afEkwFGY7E4EyHl/bAW3YlENQpKZxse/aUPOSUhD42J1rWOVEUB8g
5tKZHBR5e3MMeb3otRtezQFGlpMYoiEYb17RULfoSJZAgdhvVHkAsqDiYhvwA66Wg7Z8DhGewD+c
TsClpuoQeU5AJETdijn0RDYwfXYl9oOysrU6MbiEtm9A+RQzTphtZwac9xeKFXGB1x67F6ciJvtE
/cyP8MJhnWdPNkrje0YKxNE1/iNIFM+76C2FLSMkQEWuCNYj+KwlxYOuxiZHrXCXIZ1zfHighLKu
pG1okPEW85qtPPPVbLjOx4VQuYsKJyOdHFO36zN6mgLhZC9G7sQhUa2HkZOvXGjz8TMV86/M7W5B
zjQzzUiri7F8ZJ0BONqUT/N6KbDPguWlPdAdgywXXhEUTXmPBAqI2DzgwftxKQvfFhm9ve3rVKzq
8lOQute43dBKI7Pjq1GfsSwaVgco6HWuxaIeVpx3Ek+ZSWiHV+fskIB4xMeXw7PL54HrarVWplBN
L0a1Wbdleqm37WdOGNPyXQo7Jd0bFZtU6XVLJB4nLC/brPOWwp2NhedGa1bh6RTEfYfKNVSfdY+/
2Bat4CyI0w5EUcMKVlkx/qVkCbHFW+pZ2rsn9KSvwzoJFDapHjY3SA8udNEzG6KOGmZaSOcyrM0u
ThsuAFKzxBSG1k1yVU7qqpakPzN6guqQu1V8ZqTJvFJDa0TRQaw2325jQHWalbdKRLYjlXYTwt0v
aBRqOizvJd1OOq2rmU8gu4/Fjlv1OMbmjzmjK7WxfqN9iJkvfBYiK9rMuFJsFB2LPjlUuaOXVjte
tSVhM7j/lU6wrvsoYsPkQL/8xzQuUzqUIl06et21EcTzgirsAQQr71a2FqL21hpkxotxZpZdvD+T
nWX+omJq+JEq7GeESk3lMDrzMXA1pRmlXPZAc2QTsHHAkzbSCvFQ+RL/lHysNUeccAc0NFHNwcWc
KsQ+Kz8tTOBYOGtds3x2K9XKvO19cKicLV8Lrv6LD2KcY+EAY3pW+FjVi872YcPPDfjiL0PHRwcv
tbMVFNKbicotoWBXSVqWst+kGwmHqS1UgD8vMS45YQk1s6u1tFto6svDTtUhzCKudsqjUlDbQB/3
YzkLpKTsmydflwXvl84cp/Khx1CTFtNn0tA1HZLZ8cQqSdKq71DTr9/Zcler4vD/jDYmRznsEvNv
ICHnAEad+hWtI9DYn2IjzK629RNEOhj8NVrWpMLchX8quO7CXOuVwiZZvkrkNFhCxvkDbelvC5Cj
r88QRe9xeooqeevaSDcYvWDJa/4foevDugtvJt+R7pnFGQSRTOAbpnWZGCfnaCClD7hiRrfXra5K
uXoZzn1XjCG659PFLBXqnuUMzGVm9IFy5rvpXeGwmh8XV8nRn/yZRbnEXq5LkHoF/y/8Sm/AalwB
Rjlh7mTtvweRN+ZggLvDvOO7DRCo1KJF23+hLnIE5bgetqiO67t3zWzQ/21gm3APwGNXuChRbffA
yGfxURpPKjUIMjyQiG9yqTOBzTmOVKGm+rUd73K2KWjMXWT0wKlMdjHX34XQpZ73JdqITv2ovOTo
oWHIF/frvbfZj5EzRiOmywAL09jUTN6YehfMkBcJEys9WVCybtgLSxCTSyRmv3B52lvk2m9pMb4T
pz3D9OgxuNd5a2sG3C7XId69HrsBdlJhq2JE3nGjZuW0XHLYpCW4aGAmO1aCVi8wUdGIYmyGY7v+
0mr2uRwMkKvd+np7iypE5upxKXybbVnaG99ZnoN/A0BzA4roBdf6VcfklV2trroU0KGCJNRA5nb1
Ngbw0M7tpYOSiPzw1XlPZiVS+6BhNcOm+dRJniQfOx9A63a3sFOpwAxxEoVZ7G6FfZtAvlg2Ff9B
lGozaR/vjHuFYMj+XpaMpi+oAD5myAyo57nmRFcl7PFdaAmAw5zp32WTIu9bnx/HK+XvDuC9sdjG
Shl75kpIXt3Le6WSugZcJjP31oD7C5zeQwT9/1VPP0NlcXBcgqHONn44AhjztXwu18Dio7E2U31/
II53rLl81Ojh/qsdqG90/7171UY+5qYnt05WokGcEMNbAK68YyF9DFYX7thub8KDfjdhzaqWbyWh
uc/iydSToLSef9/m+qnH4XkkAPx5POe1JyRrqDJ+O0CF5ZlNrc2GJEgZ7LZFifnRLgvZBsOsjkDG
8/1Hl0LepkWCRg9/dO+EzbLyAKPW4KFi0ZmO+pl3ZFu4CgctNCFI238A/wsfGg1kcJHcXHlEPSTN
OKNjhvXiJS8Qpe0CWuGFjmEJdKSSNWwdMLeia8FM34rWtCQAOZnLJoefRTelIkCqZ/BdY/lz/mpV
Ob9VMf3rKSurQC6fjFRmJFmrxs9pqMwkFDIFk/wYN0p06hFhTIX8ErqD0ArWMJA3DnJRQ3OTDDMM
wFBfev4904HeSXdGN22hA0UbZTuXOry8P7zWPjnomHfPosWWli2vyOVCEcx/d4HBQKssepOb85y9
Cw3uN4L5o+7M4RYLtvZJWXu6aMnWA2EUHiKFQjdinfmKT6870y1JUsVOZ9DTqM6AVloSgfKtpsC6
in/sEpOsGrunxFEX74ETgCFWGw3V/TxKMCLeXlvNzcIvuBzmTI1EfdI6+T1BJt3mxC2B5YIOMRPa
vEwapk8v0jc10gi9hVOzt0PmEcY5EG71FMVc6QUc1L+vnBb+beH0MemErPEYAhUzL3xskXhoKZlS
0USiHzvEJ3Iq/vipLSfT+gys4nN5JfXPjNrivi/svpRy2Clqw6bvSdCvacVIjoPFQ5qBk15YMETq
5zQz4EZ1TR/ZWPBvBM3lHcWxhlxUfXsni3valoBLDe+SaCfXkq+gZU4sd+aS7kmu4eYGWTPStkXw
ygNAND1nxiuhWaOA2RigisKJKvjDj05ox7RqPxMNiCUrk4zQ/hxyEKyG9T9Og4hObmCrXGKQSlh+
Y+vuEp1+LQbYzZ1gB/0WRnfmA1cWscS2wQA8YaNDjZn6PKsEKF+pIkYh13MKStYZI+Xkc10xMLtP
7VoamdtVThzHEymTbzoSFoxCdlz0lJPDhe4K23ywsuYsgKeSCick8z35I0tamHmDmxbwgAh9wQwS
Mq18ASFZA3vZsSKmaHzrTOt3X5TTJW+h/6oYq6r4n3NvpDulkG9+Mm7OPR3Q7iK9qLJF+uFyuqc7
MQvkenrmkBdAzaJKAZ3AVZtXolHUcaYEKzZzaRciXEhqlYDAfaOBiiJy7y6Lq0oHFx0kV6HpD9T6
wcfqFrHN6Jy4r2p8Ml3uaHgr8ZoOzugFVtQN3UDTQZU5se7uhJ9jDKeSnYvVBnF+Ysk8m00Zt3gR
kPFgW1k/yo1ffh5bxZTZdkXRnQLD6iXpUJ4LYqYH9R2faB4K2+KoFMafMFDs2oWyicbOH0HCMiii
Vu4CHhlY7XPwrqSzJ3XRZbWl6v122XJKbCYf9Plfzp/J0FfHAKFx0cPqaRfUqOQsQSqU3kWPnuYO
UaDCghbWrsVzpUvzsUjFKNAG5X6uu/Pssr7E7nR2OYOaYhrlExZ/jRhgfZfbXILrLLAZv0H+j3sw
Em0y2in8JFN9NtbiYeXVEp2KjjJyzcjKyVF3Gpf3cyn0/JzBoH0BoAkkMIRQz59VF0J5+jVmI1oz
xeE9BxkdTkHDyBUSYVMfeyvHDqT58QnAmBak32nmf3ch99/w3uDbTUcnvFDyDiw3c6kmzS4I0gef
0s9o04pW60/HuiHXCAIyMM0d8CfkwPLHz/TkBTfIX88Vr7Xq8P81HwRU2c/HY0ZqSBnvykRRoX1H
J/rK+NhNugZS32HnT7xA92T1PT1SS4TpxCp2b2pb2YzMA6ISQkBXa99+hb1eM5ZnUbz/iYz5ENCw
jz7eqwDODJiXVG/gD9aSDfcc9WNmxkhlsLkzNmPxEZ66GYwzrIDJXDxkwy6SfFT9BPfI8m9nmr7g
3cbPh4IEAAUrS80ZHH5g/3LHZLfqCSQFawkLnECEahNklNrXBJGOKhApatCmNbsuPnbgqWdAuoj5
Qk9Ss00/vpYZj980ja5xe4WSu/o3KGtitAqB0h+h8Hr4WEZXVLcllijfSbV/LRmED8VisQiGwOHt
WnO+u3b/Y+U1iX6l6D6H1T6XrFGR0ySQ7Vl96DIaaYWpOE6dbWZ8WrHAJui8nHQJ49TkK5kdKCtL
5nK8c30xIcsSboNGLFscoi1iMhNkzSdyAFDtJhF/4ekrA4R98Jxavk04/FbuZ1F/wb/bcZnPBlOF
u2UuywJB1utaZM8Z+TQUJt/b0xBtnC3m5wnG/9Lb9B63cgobSzHDHVoNlf08TBFEPYPZc4XtlYzF
eJnuWnH2jget0YbIOn714p9bMNi7yaqnLumYVRVdce3cG6fzVEK9Dohqfb/C+WPsocxBiO9k2jG+
0rawLeP47YHVK/AvocFvy8Y5meLz1FdWryRGFc1y2Td9Nv/b1BTDOTDc+J+rQJJEc9j502tQLt9o
PURqhDiizZGmUXB5iFb8jbsw/7XxvAaRtyeW+DCWrpKrF/SqKBhPTzSbTgCRB1boNoWgXl4h/PL2
NjsUEDvLE47fA5qQbJcUN58vbFuSLqwaIiwbsjK0lOygibOlnIHPTASNyrBhZ6zbljEXM+ey9rXH
Sbx8O0rZPEGctPrsLiPse+HqvBMX3fDP3jmzUCbZhnjiCbceDr9p/6RGNbdi384JYgQowWA4wgFz
Gp24yq/DJIDLB6NmxAbm8d65oMKuP1hjsOTK8sDNKyvEl9jKU9EsmT4dOUe2t54qZpCd61LniNzg
C/SO09I52nQDF2TB/RMWoFA5175QgfkdW8Q4WG2aUhBvVzdKX57tTMZfh3x054qsZ8os+jBqGJWr
4PAES8HbYJ93oW/dxIRZfUGqQOntErTqXRrKWvvHqqSPwVm0TMlwb3kmIf59saE5HrADihiEJOIK
41684eNV1vNf7WibNWG+Kxi9UK751dCBcO1FsVWO6fEwE4kY0GVXofNMwhcBt0fZW3b22sPpyIbt
wAMUNUc5yqLVZ1OwOisk1YtRyYt5ymmy93ui9DHPkoPZCvvoC921oHeDbbPT+TimdyCnIxJDyaIl
vLK5fv1783h16gljbG3WbXJckbiCG6HBGGdhhx9mB3iQUwvUY8A6Ct/KABxcF/36m+4CXMpRu2kQ
1POHLEZENiMtgs7XmH96He+SC5ri3qu2xquGlLHaTKCOOCF+hEFQMnwXyFFGAd5MFDL2Czrv300x
LGZh13IdPlnzCvdVLgf0hy5/pgfn3B7b8O/pqE+vV4Ym4Bos8MmH/+ZwNAhyRMR5WNC+lYeUQ6mz
rqSnJKaaYiPrp4jVvofQMa1LGx8ns+aTyVpieOZy3RkPrigJluKpnr6J9p7myXQ3Tu4TCil0KPl5
zsZ/3xtf+Ur7FYURqcuyoq8WZR2QOdvBo6oBEtsV5m6aSwTsWVIfwyv89ybmTunG76Gy6OF3nSF8
b+mMj+DwSJpaBIcBTSacR3xzflax3uVo7wsOP9LfIGjirHBWLu1rldraPeNO/iOFtMybBmk24tnV
zzdT2GqHInD7jUbTt4+N/+bh764bkzumqqsfKsPQl+2WKq+Hrrwiv4eWJzcgqxrFsgvOxrK+Mta2
Kjip2EKodhoHDo5nc3UPPvIFQVKLrhJy5wVNabZbM1ncm1VHX+OesnjZX//kEo+YA0c2FOEckxJT
/kHBXSnDkkbeaDqpfBkSQZbanjta3kZrBhYQMUxOuYzJ6N2USOE0CYGuwH7dDaqKFPdMAcc651Gf
u2Lz+CDS12XvcS/45bZoIGR0uKF1+QZmKbVnfGceJ0kV9Jk13Hxe86PfbsmlBwIJDonJHQ67Yfbp
s2YZDd/Fkh5bNQWX4vkhY3NMPCZ1Kyyj/q756bQXt2KmTW7vVQQjRSVUcByIhWtutnns/ft/b9fG
OzUa+crOHGgG/bRZ3FnKyFxVOqvI6FRyWXhVAU48fxyw/tLKUrDHX65v7QK+yZpknjGU1e3fHvZF
yze+kElNyNcYN6R4d1zxk9t1ZSdgzdUpzzLE+T3Zzk33mf63HCQIYCZgiLsMjd66/dJuC8w+YS9O
eL3+3UgkAZ2Oh1sxSmDWlvaFF87JtPCVoPKvTmiC86gQPdXzlMRexDR+kO57GuBD1ym3COx4pGdq
rmUs5gZb+aHHdy4EQpWzaDOhJKIJHE5mZwZ0fJcnVMh5NQMmTI71oItIfcRTPdx0kzx548bUQimO
SaWluvhMERK8qvC/ZvH9rOfME+BppDfnRkCmBbzh9TiGHuX4QwlQWbDaa5cFCMbYc8unxbEHrSe3
W6F3tZql7IzSsMreyZhg9alfo49lCxgDdYEODL+49yM1Lt+UUYfHPpcso1Qd+osYJ+c/jIGD4zjl
w2fWNqI2RfTRBjlLfTM9BrigC3eOO05JqMT+htG2t4K1nMZ9vtfO94iDDjkfeifsZ1WkeQvvK4cz
Y15CcC0Jgaov+Z0C2IJFlpLH+o3nPHDX7eExFWZAnLcBHqU6Sap344k7tMT1T2qYxRbLRvqhv+fS
AD/cS4C/9Ac1/WLPE5zW8O4dcfoA7Wgw7lIviIclbtVaso2D2IP+PbBDtwRZQL62PJTipA9NZcGm
oJaNSnPa/qIdVWWNZlYg6PkSb9Gs5pMbPUDyBKWNeUtr9108rThKpFP0NL2zKEl/lBHs3FpUcNJz
ymZCXJiKFbEkEiHVVGe0m7MjF+FEBrfT9Fc3lS7Y+JlxmAXARB9bMyyDZWzOBXth4bQMGzuJqlLc
B9/N+PwdX3U5vBoMEwydE5d2PIERNTPg3DpIk57ZF5DKVlmq5tqB9SaUaQv1yTENatjO5yLPhAsq
wg9jzwLJD2a2tdgJZIEMKGIOgtO9KGDhb2H+TALAYJXB6bcYJuOWUMsr4QIKbEX4UETBmzu44QXP
w9I4vrqjdkx5K0hdCNIChPJvXmeYLAJ61AoyUT+Std51xawHO96FZZJzEZ/rbirFxPlIrmWZ0P8U
VpmhDRcmODG0hBXNqmAMtomCSpbm5jKiCHf6CLke90DBmB7Vw3d7q+AfTAEjMaqGqk2p1uWdScbC
Ol/q2UpfrnD45ery2S7MsFVIayWxJqyOqRornbshD2gvjGxAWLlHA8Qa9nW0N3cL91eZo+zFgNkE
g+7t63NUXHqYAGBXPTMpz//4J+8M8swTDbmj+RIld9/Ct6YsQcaqODbZzp0IXlq6ET4qEItHRjcy
m2n3nB7Skfs3CKNI/z6LDcXCcFkDyvioW46Xy+AJv0UI8AqF0A4s6zf70m/NfMj9XkPs3K/4Oye5
+oWtjPxNuo0k3Z+GvGgOGh9rZ1JGOeIaagFe3YpojPUjRy04JV4iLCPbH3yVSdRsonUuzGwTiFK4
GT8h8F2XvJx/gQu4L/JYJu4RlyqLH+bxKsOM0XJEaFNaYsKKYxQ8gohyscVujhFrafvwEZREhci7
TGv3FtEoVxv8W/wXGXMygz/6dr5v/07ARiLROTZAuXrjIpI81IYkbPCjde+6BysPwCjfsQ+ucpBr
qGUj9AL2yYeBU1QnuSrb0pWhECnpw+m29IulWeLlPJnB3NXJf4X4X6c52WIsq5UZHzJf3Oy1GjiR
QQQiqR6YqFPOlXeFsq9Vv8WandEgBsqHvgKHiPewtEX1pPsQ9qiykA3shdzXaS3dDeD8gs97Acdh
NR2wvpxPhPH9w8JDAcjb4Rx/SpzDJIL2nqy+YtGNzz/QY6rKKNezCgqyFY7b+xi3Thp4YCG3mBKO
PUCXqy7aL6nEzdwToYrIOrHgCk9qmkPdY9sj80O1Rkn8hEQnWYF5QBlUPwGiuGL97iJ9vyhp3dXK
wIpMsNu+aKgGE5ecNaxHC7Nzys0elxMMHCDp8vHM4AVsoEO2UMWiORnS+CLiSoBrM0FbHsmbA07i
fZ31MdRTYOf7kILVjIlB9bkHDoEx9smQ4n9CDBBUbJtdgK5JT1qvfvuykNam5F7NBHvYrjAXMCLA
3T2iU4h7iTUvU0ucGhv7hlpwqsHcY7lTPvI+673SQcxJ8DgyjOhJfTf90L4ZADNC/HCbpsT3xwtq
aT7766d6IfNfCjQ3oqxVjMDzeLxZPjbA4xCaKYbbp5Jh5Mi3Y7Xk5qJVAaImrKsWs8sWebEpoIHA
mWVL0ZseCyUAFQ1U9KPNVXmP8nxjYhiZV8aqT3BLGLVeaYgtkINcGcCoxsixl2XjUMAu7CJT2RDl
QcfBgjMhgqCwwILkvvPTt9EiYokP14sVh/cSb2rKrhbUAzXWoCpqZEppips/InxNHU94T1fINjeM
CFZPmm7yZSHFJyf5SNbdxcoEIjNaPIvVgaFEyA6TyRkzICmDVDKDF6S6bluZtev19mVBv16zNBuf
egsazWFxzaP7STeCIt994qIqSTdt31bYbKz5AaSp1KD14gGDDisqZktGjolhxeuU91nimwJqwrCY
T6nu3RX6tNYMebpXypHxjlySPRhJkOJ8aH2pB/e81aZr9mKG2oxtoQmnRfLq198ihJ7VsDH5CJy8
QImiSkEbDUyNc6Ham/xoiIYVi7mO4pQsVz/bAdFvC3axgNHljroqaJ1UNeKH6HSQ9emLnNlxkjLU
QlehZ8vDMhwoWaEUnoT+LqWBUxw9ng3QM2zRaQSqLrsLiJm/GAiA797lhtC31zhyIUSSf8Vz9W6n
XyiaV7HsQAFvmVfKJyJbjmh8xVGBw0T1iJS1OvAKhEju2/Chi0oEIfzRhHOTHWO+dKPa5JRI1cPY
hYf/q2WAKhZZ2sv8sQThSSdu+PvljXgTaLBOeH3KFSOATBrZqmSweyL/XlJFKPpZod4DiZ8YG/Xc
lH+h+wNczz3vAajz5jfWG4vnGVo2PIyqYVcfmjBwl3qDT/Yaw565MINI5Mj3BJ3f7+5THOeHkxJA
wBgAyJutC1hoDNNF4M1CIt/+97AVr7mkxWtBljf1DKV1wFirhtDG2V2nYvoGsC4oP3bBPOiiCbjH
o2jZYHbKN3KsrZmiW8z3iKoSxp0DerJ491YyeyGrfReAHKVW1iOo5fERx7zgpItJgQrSG1wzjfUI
kXSCwLpi/ht8Rtf/2KwMSADGMLcIY0BZhDZ3JxjNSr0BU3i2OIZtyuJXY8aYnba1vTgXHVFoogEr
c9hZce1H5FpFgcQZy6Y92//IqzK+k/Wm7kEkMjAmZ1zh3iem2WevVdHBEf1KuTwRFk5jkuueDJg5
XLDZRnhzLHU/GT8D6myrg7oIANc6xojAXhhL2rOyyZgWSw0qcdifmq14TNSR+66TNSSy6qHcNsDd
wOo1/oQbco2vwVIbbVUZLDwaSk4bftc8D4zGGivB4155WZfP4NbWalhpxl0eWDUuMsVoKHsUmfFt
km3zpsiuiPQ7pbDyJTj43o4HuYZqO/KDFM8GRUYudDh9dDFzqC7BhHEmdNMBLNmxCkeZjpRUrw4B
pULLN1DEBxvIf5HZXb27xK0cjpIr3Je3iei15VTcRzEf31LI5Vw1IEtpCblnudS44ge3LSyyqiYr
EUik4LcTzrBJ40R/UYciB9MgwaqfL+4T6mqotW5KHw2S9I5DCzVpSL7MM8H5VcRCXzirZ5e/Rhut
ogFRXMAqBnIZ2ys1EBslpx+SiPNOp9geN2PGvC7WzOjIrF2D1BrImlZztq5nFVrvGNVv0z2F9hLF
C8pDyVFykPWyzY/4dLn5aPtAEjwkGUeLRZs3ynh+S+mu5hAPUtyGsWQzxSxtOfKY5c5HJrGevcjk
zfXvVV4cs1xVTgwVa98yCfmqE0j8bVPhZK2PHIeiJbL5IVzo6otMd0GvnanMjfqUHRAogmN8wOiv
Wm37Qr1q0x8GyzX5WyLGW9lubSgSX2aJGU1OukwE+L/TRCjPdebHMExtzBISOCuU1DLwuxC2W8JR
b5P0X3e5IWrRTYulKLmzrHNJtrWIXp17zL0INLey3Dnr+7YEdrwpoe4/L+p4h6KkhhpF42xrjqbS
pULRCz7nr6uVhW3YDHG/eNeOdB+IKTAZJ37xNpd3qLDglJsDYjvibO3Dd3ESbCwZR71hhYZITykB
bcQjNCBswclIzfuauzosETrF/M8FIJQWgmNjkmSfVUyqLctjdzFwjbeqicDuFvo+KVkmetz2+fs6
N/yCQWOGUZxevkeZP+RKrOPt8hbS/vVZTsBrpMY21mCPBfYdYq82/RxODfFyXcxCcyluDpXRNTr7
6WWVKP6rSQJ1NmoiBKyGJpDb2MNIq1QIQ4MOkLqoOgSk7p8OYdc/DRCHgrdSTMGey2uaR7qX+0Bd
MknUExMr6WS1QUJURQXn8uSCuniSIh1TlfIJAFV8CzwVyO1mdVwXaORbYmGwfXmLDLN6jzvXF97H
2a5DzosFXlDqidqxvxj7xy0gm1tUxgesMdHrkNowZkrIuobdCoP8BVc0l28zZj/H2n+3zIgao6E8
XrHO0HoBGNg75xiN5cKrxvXNXyDx9cJFcKNEpHs1nR+bfLWDOvVyIp5Q2BSi0pJXGes+i2SRyMij
o68DDwcdV26jcOtaPVwguAlKBEQ7MMQh4A8B4GuxzomoxV7y4AdMYjceGwsmDNcyWZzp8+2B7h3O
3mYVWSd/GoF4E1H3D4+oqUnA0wAzOrMsYRpRp9hQe8CdTvAh038IwHDlQBFLKPElmJ8AM97pMCBQ
A0Gt/jfwwgwpjpv+77aD2epgEo0f+9vNJgaALJG04aHa3jhxNPbF0uwIQcU3EVzHkXBeeNth9KTo
IMfqSxXG48OOriDpALU/qaCKMBjD+5fixb1z/uwS52S4JCq+DOCWXgUh9kjoqWizgOOrhVQ3Zx9U
/rqHXomSsQxz1MFPcQos1wjr02j43PQiewqJYxNWbbwMK8auk8oSaXHogUQLT2+idDzMDBzgA61f
NiFjt9u+EhDvU5U7/ezpme0MfLiImS774mAKXHtCrt7UCf+y/qpImHBSUa+qMQWietKFElSyiByC
k7HW0uBwgvTOpN3yr76adta2+7vjQf4XK9r5k4Kt++EkIOjmaNKK8E7jbvtg4qefoLX5Wfk8yzbr
2gKq6Nxz1BhDfKHkgiT+8AncgMpat/iCi0+h80zrCp9YKFBsnYQ2sULLEzX9hmoxTYK0uoQs0w9u
cv/4VRW0zPRNb6lU8ZCuq2rOjN1B9hIRkO55TRmGvnp7rqBHs/43IdWfdDRgY9uAoJ1AYKt//m9z
el0rz/dKJ8DXoxCpVM4hyCbniBwAwRFaN/GOEgCn8zcl4Wdw+nJfKwJCpS8XN0SD4+MH1yD4IRtz
lgVPH77aYVorYJnWVo5kq8su5x9uu9keGDkE44CRasqXojNQYZjiiaM0d3PPPZ0op9egfEgB1DcY
N51Gx3enRPGLF8ea5yY6UhgLLjJlmjL+09oXzvVQqgWLtMScTDUlZ/1x7PyYp/498SoqjChQd0hw
p7ts2fv9VlPDBdGRjV4RsCudoXab93r8mjxUDMZVyodpsBVOjH3gZ1bLzMjxyMzo2y8WsKapJbhG
CJBNsjIT6eqEKrpvhYiqnK6njSOPoh6yE362c6WqrAeV7X6EVwpIg9/4MsOUcCE/9ytK60HBYN72
jmhsD15FbwLTZ4Mcx9ILDSDQ6JbdRsszSJFl8Y9QNWuTL1azmrivP6S5etW08a1sHZvuaAg9zsgF
y1UxmKuhLy8fOixNLYnHVQrYGWQWkRXOSnku1zCoeAWaqqByGHVf5dh3sIbfR7d4oq180LO8IVvD
weHYGyWPi7eiKrFQylKnTAOwKZ/OHY/xSX0HeE0D41JU30woURmQtj0B7g8FNySIckRfFncdcfWX
GE5COuEerT7BnDmMwpUyYir24SoGvkgypro5FU+7/tMqW3AkRVtXrw2N884tqSZ984/r6ZPRlbk1
T++epDJMisKAhIqxSqHxXofosZvfmk3TlG6dAw7Ht/Qmt5nTcc/pzu0qkh22Mc3WfM23GXssCZvG
wwjPLFq5HglQijZGjI7vFSTFSNc47lPHMwt2U0W4ZY44is0MQKncPk0TbZdZZX1qsvd1QJWad1Tp
flipsy/GeUjtJzLODBeSGFG7e/RBJzUswHI/WQs793Ud0lFm65AEMkHSHOIPyrWounObYXQVWblE
KVA/LxDZa8zO+K3RQaCZ/079WJgaGHRbk/NBq2wtJWZaMnI2JQ9M8rtpKLokAVjAG4q3cghEEj/E
BMC58UFF/3PKXwiT2S5w9GT24us7Ww2Up7DLdH3jTpB6HPIuIe9VE9bV7trb9ahZeXOzKwU6nDDX
SFCqDvpXqucvD8xz5wmZIN0/WqKRlMxkG8WdLIFfheqdRMUlr6Xi7uKaw74umEYs2PEsKc8EEPBU
3MVUjYqkf6vJTzOGr5Cb6HTxtNBMX3+qRRtlHLCBuMn5np9PRM8k9BVMjEIDzGM1TSVazaabOIaR
JpaBOZYIHQqvM4HcnFuyY8VEorFguFhs3XSOK7CvTkY+PQdx39bpa2Ct07DDvadVdwwBGJma0ulB
Jq6hn1psjb9iU3paTVp6Hexzk4JGXkGAH2Tz2YsKoQkdugPNXzQk8vxmJxT4cElI+u7rXXL+EDfW
ZjXdd69Jr8gAu+A2XFJ0OgowrpzcWef7nHEPbM69q+K4D+Vjg53PCkO0xiGI0XKz0H0n3e5wLsK2
KT+0FLDzJCLcUgPJTKTLMpxgGSy89sYtOLub+qOH71Hsy1XwjEJJMkMEW0ezt2aF62FrVpKWvKOj
01YvTInr4LX4etzROKiPJtJrPVFatYzbuylm4lCwE7bMHPIQRNBq2FBsCiaL+mxYL9Ok2cbnBC8C
irE0D3O4NKMFd6pbfXJjAxY3M1HCUFl3Wmj2uGAeL+kWNZ5UiAhe52tehhK4KX+YoFGVGaW/cvMs
iS/zylfomrv5ITm6nTA3RxV/ie671V9Xciiv3GTFgTl9VFavAhS1TV9rkAoh2Noof9heFNo+C3lm
VeiZJ3HS/w6ny/k5/+gPxgue5t64q3BVcuuayIudwmMEY2H/v1oej2iUmqmFMZ0oVrD8MysmtLHI
rTY9osNWHBtYsfg22qMA8vsF9xu7XyGc8hb2d+a6kIQGE8rZZK2IFY8chy/N9BNsTrdVBHJmXnlq
FBsn98sb3bjfTUSuaVMfKeRIeIlq8B8q6aYNPDYfRrAqjcIMpWSKskB6vj8ycWZRgwc1u7/Y6flR
raWx57NDyJPqMS+A3CVLA+nVLgAodLTw4kX0G+9qdAqRNvhIWtwrCclzHw6Ev5+TKdet/jxVQ4Eu
KjjhYSXBj+bMNnxHZPfJ0tlts3QIsy5AysNGhsy1JevmHCbsUvTgfPGUIR5TVo4qUIaNwZFPtiSM
MbUTOPfZLwkd3/N34zhc//QqK5M7eS3xWTKxuGOSJKEPtQK6HJQhQfrJpHi8DCvRVXC+G/0MS2VF
KaIABxvEJsmsfytjc1xGRRyp1PFpFl7IxphFnIQoLowovW9RhLAnL4ospmY/KVoztKZT2qoVPd6m
e3sepkUb8QH/iSysIK3GQLnAEskPRTHANaXZAv4lgnhK6gi5sVEzJXwjffIzOwzHPMOb3fHEkuPV
+BzBd8cjhr8TnQfDXzginUpJvkWH3Ju8GFe7/v1XTIbnXwMJpl9FkCF6fZDJ8NeM10pOEpzY/HGZ
AITHlpxDBjW2KIQX4rPU/2EgFfQ4kDsUoQEltRSPLiX0e8KPh9WPkIg9bPqOnf5cc5R1S74kG2VV
lQ8QS68X3TCNiAeZC6Kom5/MqHHlHF+1gi4gZnHhZKo0P8lw26Aa7+tFxqb12mLClZlXQG/1s1cM
qp5qQtmUHZuPC7ebcuhE4WbQAEttRtksF1r+flGR5+i95pp0TF6I1q7k52dTD53OoQPfbONr8FTP
SR1JmLrDAIIgRxKrZPro/5UuvTWHsj45P9FoG3gQ6npCLXRcHbAYf+NsvUUx4jnxQmfxZ4ldgERp
vTijWgTw8yxspt5TnPoyZyJmpu4hXad3axpXgcEd9R3OgABLEK34Z64mj86RMbwyCdX/zU/mJUH2
G8kdeCvgwuLjZMsBEc7XEYKu7Um0FwGvockQvebuc4187HJxvngSP6JnnZjkmXnkI7W4XUxDdAgz
lLc+0CqNGID8xhBPH/JXfj3Wt2TdRxrBglSD9+l1k3Zj8ymub3NQBFS7ou5738lcmAMu2XWrkKui
FE4rbHsCcD9zBvObq9/f2qrFwwSBH5CX9NU5aC3TDNoDSQmyc+uw8LryDbBhWIY+y1pAppNr1/6f
aZwmFJ7pEBFR6V7wBTTnqKEwiEEgwhGfH2Rar2HYaMzYF1SG7XPALUWE8RqrmhLnIFju1h57EulF
xZTt6aCa4RokwgapyHmY+ZaiqhY0T9orzsJwhd/a82497TGey1uB1PF+vrIMdUoe7Nj1XxDo2GBa
6JsG4LFAviuDTCSihswpNSu9aPbXTwDxkyEF2jXsQpfqxBikDjqotw8P2wr4afIqfW7fQH4J7t2p
88CXiJW+h2q2S0wcbgW6GEpw8TQwYtlSramVHQESOif29LloNT/g1llHNZBbGO9I9tLqlpWkSuYO
5g/c1YkvZxGZGpVEWd/H8zgRHK5aaL08JI4t0Cyv5OP8bpmgpeokSelgpYPCvsJD2+PeCEjlmVMa
XSTv0esUn/R47Lw4bV5dY3z6LSEPiQDhT6FeSCa+6RIvMK7oa5Zm7iU0mJVxJY+sESMiueHVda/w
6VG6Rgxr8w0Qj13IeI5lxBCqJCFtfGCWvacjqdkVg0rydrCKFhDFOADiKjY2dS6AJLqsWki4yhMY
aQrDFgkRmw44hLHqSqEELqynuB/I6FPJPsWpZUVoZFTdlLXqouFC/jx1VvOx1GU+W5VYURmLUZvc
Bl6h6xlDEgGQgUkpDeYbh/iNo0QpGWrZ+K84cN0dcqIFb9KYLmfhr4tT+cGX7ddzyqW6bNfwVMe/
3as26DHW1sTIliClwpE0tYr4+PYIswK8VwoCoXlq3KwkG0r6NnRgDOEqA4pcAouARVmvcgVOCHKH
gotYiLXVR8YZML+kN/p7RWK5sJfhQnTfaaiWr/VZvhQ8wWcvvopOgcPA0hzYE7KhZEr4Vlf/6+md
oI9ziFtd79cMTT+pjdqeR2IG2eT4MfPuvrpd9SHjkyXxdEqQUHA5dqlxPe+otiJY1sNjvUSkSvbj
obyTW/qjvZldiSYwsO4qoNpQXFZ4GtZIpbTSlVeLqt6K8hxhvpwjBSDNP/cxseUTBCwNaunrKlyK
RvPS7GHP9rAhUVMN3BEDXwYcjgPwDjTMzlk0kFabHjrJ1IQSLz1G3J7e/AmtxCrYuC4huRaBgrxY
3kWuDoNZaGdWca7y1xPGqBTHyc8W93qe5X8Xv7oMogkXFj4kjCp5RZuoJmjt1xEFqEOaR0/m5TCc
kyDt/ChWAOOUB6ShjObsfvvSx4lYgdHWPRSGL3pBwGBcESz4a63DzHV40t1B5eGgu0xZ4omoC2mD
DH2dg/IQ6i6APIV3HR7HkvSq3eSfK9LyVtdXosuJRzYGbutG91jdn0fP6Trb74ml1xrhf/y/reUf
2hYGUpYNxBQ4FT/75Y1PP97Tza+5jwtw8fgtxXBUKp5fbuUdHp5Gbs0szDjDEW/5eH2uWPNmmjer
yIhbS6F8kWn63ahYJk9cVyouiw6cfO82/Mb/pgEWrTloWi1VfrkuYC4Pg2Kf+x6n6/cX+9CcA7fP
sEYJdUnETCjd02OVXRf9/ZJ77SuKayM4e0N9TJJfBP65AUXtGz2NDYi1REvqMloYXTZeyHd85kxG
Iqm2mc/cWVUuG+0b1si663L+gK9FLl+Gwy2jcNvAfUz0F8LDns/PEUo2XJRH3D7Do0EEeWYTtsBq
Z0RBzX+Gnu/XnN+oZ8Q/bXiDFV9vJfaOERpqvLOG+1jzsMlXFPztQ01fVc0O4vFi7PibYy3W56MS
Eis/nrnTVmsqPqUBAIibglVirlii5m+Ax2Lzn0fz8UAFfMdgUFBjfOktGxhgKYdZ21uW1wG9WNie
CF1f6pAl54Z1B3rWllc+yP+8rtpo8IUT9lajvryuedkKnF48godfi0aEj/U6KyiFS0UFvnFY6S5L
V+O+ZVvIKtCNXbZVxdNSVcVfrQp8tG+0nq+ChakcYgkYXgbDOvOIlsALRtfmBI2r87/PqZVD5Ffm
B+LrGL7i2JTCMBIO1TgKWiJNubsfqxt3QiV9RK5qx1+e53pv/O2wlIQc8T37Wv6LS7vZjqB6+L1I
KVX0hH0ByvwafpbEpk0QR93Y7a0U1I8aeFeh5Na0QdQ8JWv8RYTaD3ouTibmAyQGPanp+l1NDOiU
Qpz8n0JTdRjvL40xXRFC3zP94ssrdogkXxMcXc09KfQhUZkt95OsVvmm5dtXCRGYBovCkoPaiUjL
Ryp/0gNRplwd3MXgVqFwvh1jPQ9JoJiJT1IbH9XBe4Cq4s9nDXOUGpmV98x041vu0UQ39R5eHoGC
gWdIBfKp/9u4HaoHdC7VoS26DUIGf6Qdi0ERCbiQTMGygyaBZZa8Sb1NdqaIYIu/KJTV1hxMI64x
DMoZQs++kOMnFbX9ouTw+Fjuo24/sx8lZvgzNJ2RvSwaxOrUyydR1xcyq51as6BO6T5NzW9vXq32
ZQ1SZ+io6uwB3vqq+opkyEbNktMeOTAiImJ7psN9UZct0hcjALUksuADDFMDUATlrFnTNz/XvoH0
f0kZpO6SEKPomDI6cIgvT00Nq1LNQHdNGILqQb+aKFUrjKltXVhTJ2D5ePkn4iKMiz/5/XSVtyEM
eDoHq+yqA1aX254ulWgmI5JEZwh+wk5WUeqHGx6yCfrv1YusCDBM2XTP0Kd9y3si2jJmG8gfNJw1
oE/CY3OGEchrZj/nWMf7CQBbBTfT2Dx/esAubUFsmk55bGbnePIQo1nJPD5emL4nGkbZp8NoPD4a
GSrtJ7n/TbQtjUY1ZDR3Bo9vt+1HpeqAwnjctUOGcyL/FEnQeVJtGfEEp5xi+84CCbDlkNhjctzC
B4WPNqVk5+E5qNVWEWJhJ1sp0Sw8OH+dj5APGQB8dSSf9M7GG0I8x9COLVb4Cr01aufZH3+Et+wY
l2kCQgfvu+Ue0cX6VQco4tOePOmvM1mWrGkqrXN3g39rh8fnfGmBTqG59gy35EHgJK3JFXe+sUJp
4MQ/MLTbzVqXCFytpPvfrGl/WBTpJ6Y+Gw6yiE5wQvcK/dT2/fP3K5k80+LzHM1jC1Rcd5MsNUCg
SBlpJLqHBFJa26dWLXSeAHWlnhawFZvvaMtj1BpStzo3DiNp8d8GTwM0YuDpXsGl8iwVi3DSe7Ji
pdf3QJECw4L52PWV2XjVTzhiZfDrJXJleok7xyNhgmfeNef7k4l86Ik2qEl4fYxA/HfvDHI1gcIa
keW6W2+VjuyOmLElPQUlqYEt5KZb3G+t77uW99+Vu9tgX7/COjOsaF2BTtieNfiy1JvggfM48qi5
HE9Iix1TnB7AjmPh+VOeP1yD87EcZIO9sp/xPDMYtzV8LdbPJAPIw5mTo+TP90R1KuinCC9HVO4e
+yl3Z9k+W0qim4LKzR07Zz9++DkR4p9xpv56tUxX+MYUgaMyZJO8826H10EazvTFJe+96oyG/U7o
OihUQT/PpTlV6TfFmnv7Giwu5ADxejJBdPO77U23iRXIIXnVUnKgRQUimZmlEJY6K4F2gi7VNQlV
W0yFhJZY4RhFUwqnUdSh7/OMiWoROOoFhRTkkKpT2XUBZJwQfre3iHSNNK1j5m58orKQjcZHmZ2t
+pUUlX417skJNWu30HhrofSVkBw2KznVl0PMagZDLcsG3PcFZa7QajFcCUiwUVU+uDrrQhNfCvIM
+zPyy31R5wUxQCKf9HYPW85fhpEpzK035Fd/G6xWMWRM/VH38Vo06wC1TrO6T9tWw4ON00jemrL9
VLMXbGrmj2qi8z6MjOz/KZ4FG63XRbva7F1fjue8rJLaMX1K7gdmmV1if/G1BcRMu1Pum8BJBhkU
Jo22la1PfbEx3IJr0AFKcw3zOZdIkFDwgfLbDadArTgG3I3CgKZkmbAoKYxUS7+GLvNXN0H+m0MK
dTZ+bXEiGFKDgwatFlZMLDq3oPMFRiaLjLO6+WiMXmvu6HJkhCXnJkZxxN1rfCK7n+2usCMPVeQT
WZEQCcV70VMDxqlLf0mQoDKONf5AAUdo6wrSI4XreOjoMyEFk/AqFm1u/Ac7xEJuzIPVS/KnSMxX
kH3Lw0IZKBPL2JEmjBbLRa57g+Oc/+XQvZ6ayc/ePxE2lGaTdZ9gkSQjmj8NLX6bOWzLwoA2xvUq
9s6fol501vrc4E4oG8JRoc0hN1f10Z7q56k6Do5o7/Oe1thiSnQsS0V+4H1MaCmEIPptubNj0B3u
d77ctNUNWsH4qVK6xe6vW1KiErgsO++2OUxrfvV6K4vtGLwkwT03k1R18r0qRkrjtrqQROLNiKWU
D+54xlHOHzu8jVdIG4llr8fllB3Q6SD8r+41hS8YC+U2oV9zz9Oy3G91OP/R2zihc8uFQFOgvNFD
RQUd5LGNSnhgyftwJqGi/XDTsVLyqlOe7WbLK9pCioJsMTWWU9fgLgq8Nhwzz0IMvZhgQgloPOmY
Hp2lkkst+A9vvH8Bi5CaEpnyQhr/5YKQRqZp8SXO2QkM7Nt032wQC5kpn0Mu5lVjDw+VFbDtNwqQ
jfzpanLJpY1IxMerV6FhnH89g+t9UV9f912kXJO/tWDsaM9ep9xksM1EkpYUmYxQNIZS4A3UAYDZ
Qq056oqze7PAvhc270cm8TXUg4vMo/M5Lwb+Z15uDK0s4efdcy8fubLUZXiT+WEKVA5gCkZPg7f3
+iMm1kmy/QYy+THsEpyEqoEKWYKjiD6oPA33CvG4MgtNKR/QaZLxppB9ldSRrP2kNm790F88ZRb2
H33hlnwN98rahQBHwTLKJ2eddUYdHvdFgDqO84Hy4+xUu5rPM0p5QGNQBPdTFM3uEGa5EFuWQUUt
KwtyVMuwHJp3YcbHoPVbzdNGCoTWTUAX9+XB5ZfKER1rBEF4tezgsbKyyJn+W0JogV+Ra8afS+Ot
n+ZK8mXKX5sUw86uoaX6D4sgBI4PuwPFMfzKHsqcJJyKtX4Y/WV7hjaC+uoN4+XrjshpAPL3lH6I
eO9JcVCMBTzsdjaHR+DHx0qcDGOl0lktxf4ZATC66hyavU8/oCKmpJTbPfXOMCy79kQugarQBnKM
7uNLk/SH5uYRZtG/HKWvw1VRGwHZlUCEkFNM5z123SXajhydy+kNgtBnly2o/INTALW2hKQWuZhY
JdMYqS9tmZUvGgBhP+eDabXSjTu7EksH40/O+VVTX++zjfUFJMaBuib0V9mJIoQMxG+sMkRrGvNU
kYiz7MnyAelb9jaEa7dOCmJtNhH8yQp8xxrYLOZsKhd3fdzeeVuJvI7WK3lZhTrtK1dC7THpG+aI
Z8ecJzUCcHKgQac0ztS9nnxCure2uw7DJeASJltYFO+UUCSprtuqL7IeXqkNRN2WO+YkGwSBdDsB
0cCpo/w6rxtXXn1TSqgMzu9I3Onwv8Jz4Ip278S15REaMHRX9SaCJzIjcxkjKq2XkzjSNo4prAF8
9x+azfrKdQp38oBmX5VWkds/mADED0ZAhpJNaYD8BI9FHJo3Gt8YG6RJvQOIhYXzEenWQTiyMHRW
0tPjZzSF8WEuDZIRmcPxJUYyCQMCgBSqlndM1zj/sUaufvGFpoRFLbnp9yFet11phlIreHq7dh8P
ccS7/pxUHvtXIcIcOiYIV6uvRJ7bJnX4+paCkvOllGoeJ2YKr3HHw/2NUW3j0SasEcoDlhGMNBJ2
2uk9KMu8O1i15Ha4dK21KW/l7u7n8/Spc3dywKr+uHAgOBJHp2U3KmXPUs9wMsvDy4BX2T3rgi4g
Jbt6aPj2dTCVRid0gaxZ6iFb6O0m8FgYmitRDlFZSFa4O/ZhQ+WhILzdo59Ko9lksShe4tW0tggZ
qAOQVF3ZTr23vO7nbMtJ4tJiUYzpIEzQX0UZjGaRk/4yYQCq1wA4X2sh4snblsbSCi6uZ7UFdW7i
GRHrEPRJ0xOm/oh2UWp02+LFyt8kk5OkTgLVmF5aOrRIRZd0y1PKrpsPcLR93nxshVLRhyU6VSEF
IOt7jp4gEcnLTOMWlootV3F6cC4vnhYxzpsj+6m0wrGLdyYPVR0xy5zqVZJYNz2tLkSIQKuDtjzd
/DRwFkw10XcUnEhuvbTcSGHdcWIA5rNKBvM8ppMUeIv3v+lD5mdr04YqnXLObBC7300UFDEk6dlJ
C6SlApkOZobuUHlDzIRiMKpR7WS+K8qwtvtmyKgF6Ysdnhfa7/b9Y/KZ8N9NmXSeltHI0ie3OJM1
tjJlENJ/leYgsm6ZG1PpIFVO5kcFZn8GlP9qKbaPMDXr5r1gdrJNU5uUncQaCghQmYrEgyALvZcs
wS/MkhHltAUsloHa4gWrT/ZePYWxzWBVeRBcpB6txFXRlwrXZdaCyDuoVqiWVtDOX4EsGSNfMxl1
LGSRbjlaNyes3iTmDw/9KtvnLZ2Jgz/U9KvcHHlUUjyWNjaKFUJkmKVhCZDDB1ggAETzH4AjsMfe
k1NHY9ySO5VP02qjONHiG4wDx0vMH2ktN64HcDKkdGxtJw5qvZVn/YbUAilr92+xB6lqVGM63mT0
SIKMl9Wcqh1usZ1D6WlL3kVV/w2RoCcsyaynLOgIkwFSO5xHQtQWAw8NWyJGRuJ6TteoF0xOBlIK
1TlB3aZxRpDK45lVuLNC/Do0hCsYUPk8Gj35ur5t+/ZfBorIDtcKJ5EBVGVJlhJeeOnvGG2rNkHq
DRrJPHtj3TvlkkDmZYiAGa0G0PzGCje71k1JFEJsz9y6w7yuEwXEVtZ5X2i6pA5pDA8vrB+2FLjn
4SJ6JdgJ73quMrOP0mASnHma2hqGrSYdYc7B74D1z+1jT0rdRRpgVyiIZOF4UmuIEuvBxfGKjMiR
a/8VMirTzGVv03E6peCpjsIT/u+i9YwfnyjGQ7QZalA3iie6nNugoA1V7VgUevEbiMJH4ODiji9K
tYt2RMxeswU/uwVjkH7MUq1tkeuONwJ8K2f0EasVoa9leKYD6pjlwPN7H7m3lag2M3smYnnDrMID
osqGj75cDOc1WBUevWillMjMQyVhkEI+dTu37Jvk0daOcs1F8XPE0FXobWhCV0tegfO8TtuwhdQT
9UfuT8rnI2fm1PUt/Uj12GDhvf0AeUpX9fe+rjSBZ41d5WRUofg8n63vuQ2AccQzvi3+kY8maAtT
+AeksxqCbXUvgkaKAGOqw3B4mVdElBEo04TemgqOpuMDGW8UJndoFHIKpG22rOIeyKY2WsdB5cOX
/oVMaRVOeaj7958VNu3rcjO+blEi6wZB9z74yPTx3U6i27yq7om8UMBohmlPJ+39jkrBKkeUEn5R
crpvovbIrcMhBrPcVUQ5SxcQZn3IEKr1mJCLmASv8RTZ4PuljuMlVDXTt5nL10wU1nwdMbV1T8t9
5hNcdxi+X53roLnK+yzYP3Zdwh0XI7UqMTIbIEbWki6QXLgbWZWBhBfJGKOteK4Zx5EuPAMk2rO5
+X2HdcPDWxd2FBXegdLz5Uw1NZARlkT5bXp3aYMqBaJdQ/O8jOIltNB6sis+wNGmvN+croR+uqTZ
puLspxEx3FXYJpCE5nE8pGVNI1qlC+TOOR5GJnszDziWS2MmunsuAK4oe7aSw6oqLjAArefCmY1P
8F/VoSt+ltEsH0X97RiTnSH9H9Mtl6qWGJ4M6qrllxUcQl83UTRu++nbfJiw5IPVAL7ZeIhtzNxc
Zq1+NZbUBpiozWrK0ClCbilhrLhywgkVXoJ4F5ng414RjDFO6DVGJoA/yBGwYTDqTRGPjISkLVFD
owWl+rus0YHmTWE4Y11D9jY6NaCedOFSnee+Nu6ylIFKaBYiQvgjO2IrKTOlvrYYKvPbaALzKJq5
fK5TeJqavsSXwhiGK2FuWGt1aGP/Sq9EJDxyOHUCxdNxIR+hBHWuy8+rQ6IH+fosGkWj7HRVCx0O
M7Qfpcq4ccMyJOWxiMHSIKjSCTjGg+bZAEeqdzIwn4lowvGqyJxOqfTa4Pf2fY8Qzej0vMYKoEej
NsadW2JbTWAbW903mKcwKCPYFgUXPM51OcoAm2kLHrtWjBmNK18lQZ7iPJUacCnhYB74isbEaacG
QqFo3NRdXUkuDYkavUJi4DOc3WHxLwePIHZYbTefdIr0NF+3Z3IzTdRmM1mHuLUARL0cSZSgTfyl
3xjyb5pcmht4AUbGewMlC0r4WT4ZwQZ5khjFHfwltWxI7H06jM/Anbbak/QW21INIXzBGnbgT3EB
V0RtBGiQl63qQLVly10/EjaFLjftKGGs+zeZRizlKB/vQg4V+f1Zfa/zuokLzi64ExIO99l1xBRy
Z+3YYt34AVyOvtCylQyitkp3T2ZXlxs5bH3BHmlrDM1Mh6DAdoqe5DynPS+GtkuRtytl0vpq3sg5
ciBhLA++CaB6TAhN/Y8RC1RKYJqLwbRYs9Ro4hmUIprsAX64JV6Uxwoihuc8zY1LKg1VmcnfDRNH
QopFkZbDYXlfg8srqgSLZOvcciBMCzvw311SqOv+I3QEsSdHYb3GdCNlIdBxsV37K0nYJeGYUd6I
tJDwN8GwrJ6nNxFGV/5cu3yeiveYZ3jSzYelRn883VSGHjdWbU/kTSO/FpmrqOptHsXl0sdmHoN0
Rwcfr+OipLWB8NMq0zR5i5gu9PkhWKrZzjwQuriG0Oqsgf/TbbeJKBVybyWpgH7pLPsHKx9zW3PU
qINFE5MTWVDEczhNj3zSHbAJ2CCbAHd9lLa6NuUa/ykQEH8ZUFkVdIbgzdej1yBuFtHOIt9gUtf9
E25Oll8V6F52wVUX7Y3fQElDRG2xrA1tNf6Z13dFLHlrT4ymDBPT0cyj0IvVUTjSLncvK3dBWaWH
ByIJCNzLSvF7IPr27iqnN7gw6/AMAc3Kx7Buu7kN9sNskR8ky+NTAxCyQOKpgaASAatBcSwIroKa
rgmIeY40UErPmdWo9gOtOpumSUbdRpG26dmhcz+yLmekxAT6SJ4D0OrSMtTceLG/rv8nNhArR5yF
ekiyt97Xdce4hWRxwQDLB04qgjpk0LKTD/2Fgx5nqyiyz3N0raA/1F8KRskxUEMi5MBtqiLi4rKO
iBF5AStnat6zXpIbNvBwTxP+MjnOp/P58LsFlhTUrbs2EkmSmvgdLbxMFgpT9bXcpsbAhw/BmPy7
qE4TI96gVpjcXgU6gsnpyB7ioWZ2xVcBlTlUE2R0WIMgE615Yy8gd7eQ5SA0OqN2ELvBiS4gDh7H
YZ4cjKI2la0u6xrItjjjBHdH/taHeCOuUfHuS1edgeOfM3USPj/7d4ILcsoRMYRYoFPSaHL2XSqH
MtToBj4aFW1ifaWefKXULzuPUjCUJ6yccwRuTQn1+WBLWi6mke24AnnG3IVhy1clBH+ZaFbE2WpN
sYn3CKcOAF2tAjZnEtxleqvXqFzzLhAVxTtGvwPRnhVgRDk6vU2CaL/NyNDGwX1PixSYJE/QPcdi
v654y/hKgEDmx56rRlhUaavO9s6kmT+pzAQcMDfNcEQUmaRkHphSjwo5DboiTS4l7ONdy6sA9T2N
fGWspFoc78IVw/mscZ5PTfJ2rXuuQJAAG2ItAUUD68tjS9ks9owwBtFXZHXw3SDdETgYrTboeAPv
ClUar+sKE5VCc2SzMCzCL0wXt5GfAIYPHoNp3TnYES9sDOqC87mmRgY0hgh871e3kjD5KUP8jfNm
9vYmUhHkVH3h/DWypCzG7Kn3SmY+fxF37YByll7OX6Ju/O7jq92Mw1DmtBhmt2YpzIg/7RrqUANB
e6G1t4tRlo+la1GpDvi+nzez5Q2t81f+ei9btsLvxzbZZHSwsnIf1HzbFsC9LEBALmoRf3de8IPk
YOEINZyqKsoiAyDjz5yX9pdDrYDL+Zmg/Tz/qhTi5nakFt3atFx/RBIi4NyAeJDPmNj6lJ+T45d8
9vl0OlrEXKiEfp66dm1C/jkjo+pNs9vEBG0VChsPWHUw7n68mVQibW3tpfinPl0DlCEibVMzUW5r
WoB0ywff7aZAdVZAR3U0zbJjAegcUN3Jm0vAmdUunQZLY1y0J4kaQGRDGLfJ08NHpJzszapm4yKm
BLKIKbQ/BsQiylIhnrYhwQ6qs1eAUosgt+/8XEPKF3sm/qLRxh8X9MKQAdDMgtPaUaDFw87jS6RL
Y0YC4pfpjDUkFXv2gQCxG+JDIaK50mTeQPPjZOZVeBDICAsG+4wkLUqa8X1np2zm0dkhVCtqH4ju
3DX9PXKLDTbHcr+AcKH5+A3e401TIE9ZMaQf5QX9jayNK+YPW0UpppKfcZ10uERzvVnS5no6asgl
re5mr6QtRXiqtHnpO+2Fz5KE6aF97LQAIluGzmjntYwYQBP8a+eCtnHvxbAYMPNuduRt+ODW/y7u
+drr3iTypELSDTPLrK2mfvwkWhj/sM2FprnHihJW9sogTv+6GOe1qJxYlMVkw1W1huDmOgPjMlF2
UJDMexqmshCzCyBls6Fa+vtXQ6ZC1kT/i+Ye/ylXNmlDlV1ph6wpHc6t3joA0Zbg5BwHPMFkINv1
Q7fcWT5mLR65NstpLA5Crdou9xbOoHN8XzVGadkcJKqYrSyKquKT2X9YS1gWynLgvWj/Qh0azckx
ooK1TMYf/16fJVlg0fSB77Ah0sFvnPJXL5TdHGDeDLdXkwDNtPEHX5putpE8z8QGoZYwwWuuKmms
EzJjH/rbXkAWXG//T+c8x4lxuSgNRMiQ+rYn2I9daskEpBPMPzr/ONWpybATMgxHp+JnL/SjnILy
/8nOBNqotCSJoRYLl29+UDcVQcWag4KGY5S8OcuL5qugYICi9H9rD3JgJswH/iF+iW1wBCxG0Oq2
56rOtEnmnEMWAab7BwvlW+4kjAauj6NoVUsvACz2tfhRaJxr4oBvDHanRo1OrYRlkhLJI4oaYoF7
aB5GJSRQs0uTz+C8YKcqFrujqmvJ/GUCOWVbXKNbJAMMQtBjPxrSUxWm7joX21Cy55/uFCpynbxf
Wryigu25kpDOgrNT5t5DlN4+HwL4tasBlGoKlvfAhRndihtUYqphxXctnmO8DpQuF1VNP7nmpGzJ
D9H2OyIzDGRqrwG8jaO7Xf3tQt6jpj2pOJNyMaaTjQ3h3wWcS0Lg4Pou6CT3/aED93pfeoTlhgAF
t9kV5ASs/jaFg2Rys3TQ8o5UIlHMF/q/dzehbUvBAWNHzyp40YFf1PR6nOi1cMTdgIqZMpYqzO6V
0ShsF7j6t4OdueiUdyjZjsdwt8NwFR2ajlI1Z0jBHOgNeaMp6dtt4Gz45UBPocWttzec0kLfQTk7
Rc5eaPLKf7yjoCiLHQuCaLLXXMY/qGDPKzBtC5E+HmrVIqNAfoHHAS7ZeK7NXKOq4aUXncMcNDNQ
NeB+1XtByC7KLK/kbSJI/nLjmU/pSJopFAuH504PRzGQ4Ljvg3zPxwf7l3s6oJHq275NM5zDW0Yl
RiUUybY08knXjVudETJ4AH5SvqQ6gHXkXnhCIoT3Y7cLc9s2abRI24qWyilQnDO4dAI7P3YQQE+o
cOjyzJdQLFlM+vV/fnYo9jCHjjKQIij6Akb8ZCtDGyX/nYyU+BYJsFdCLyLA6w8PuScFSwJ1nAx/
qQBsf3JVTPRw43kFF4pvk6CtN4QXzJE7gvDk1dJ9GMaEOM3nXsd2UOCfbdCzOvDMhw6AEMJ959uF
sw/s/1tRiGdvRjifO9hyCO/jRQMwi9ZN96Unm+H4gjGDDCCGx5Q+l7KcMdrqTPOic1QCKLzvUSWS
+FA3cIIRL/rh7VRBA+uvLs0O2tIXXyCL3nhuIQdBWwyY80tiI4ZOPryToCGLFenkE1L18/ipcORD
JpZYdUukvi9xTj+igDvCY3RU3JgdZ6Z8sIwh3Kq8iAG+5yK+/qVsbIkHhIU9SRmR1P7UZwxNoCSw
EG7NhY32DbB1BTXi1lMh8M33AI2SfuS7tRrdM6AwYP+8qM9SJnrnjfu0hQHtEupRbgCbQ9ypQaZF
BeNABnKwh07ffpH2Ivrjbg6N5zBiIJm2psZnA2Ob6ESetVtuXn0E5lCEbwLdAPPEyZxZSuhgbNU/
Pm2lY0U26XnY26xMbE8b7hdvdEMThU0nq8RUyIjUuBD1gphn2O+S8BHJx+e04coVf9DxufKEIqKv
s+RBkK9pHd2l82VanEVH4zDR65JnRIESsq2rjkbkEttzpv88IocpNn48iCVa9DFnQvjWKbAsX4e0
/eJwjBfHiBOh45bEmU2H7IUgb15FtS0Y1GVfmrsBOyyXyodSBDaBfqgIN2iPuYVKwSPSx4qpysjy
eyjVxEOmcFwTTjkxtmGyY8+WmtsXff6ruzmrzZfn3Wkly1NDOWmisuQWvDpAZYjzUDHf8aqGIL/N
7yXCsIH6iFxCTUWBD6EYSqucoHqHGblxZhxiPmB8jwwwk7fle9mtbyZyLP2spUYuRwuUT2ZuZaK0
3CFHwXJVkhTG1Aj3n4aU5z+cjFbvr3WuRUyTapMVCOd+WaFjPYgdJmhBSJVt8JdIvU/yPy6lbpOb
n5xUuTB+PLi/9pPF1lFNgQaZ+FMW4IDUbTqZMAZzgB9C3+2ASeeDCQ+vhCneQJ2uS5DdyDyWyZs5
wJ8Tpf4e5oxhX+mTuUjOsanGZd9z2+P4QQWgz0zEhI9x0TIDq1WxXr0M5YCWVGlb+Naaj8Rupxyb
xONRfrmd05SQFhNOALURiRyMWdayC40HDZoYwV5tlnX5GI7FslzPOnkoEmu0QRwkZF/BMotOCigM
+VeiINV4HxOQZaOfahDdd6IA/oRUKqxxUB3BRwu+pASgCw/4FfEnD8AxqoARd1QPm1ihDmVScCNO
/2LID/oaLUZx7v4QniMX4scxJEKtzCvlVChoLDGwjLXpDIMQ7m9SIsv0RKWgLtN7MjApQRVeIplY
/3e97ZQNQ4dp/1Bbmy6h3Vg2+C15eh/XMRvbVpibwNUDhNKatLCRhbL0F+SOxzP1FHgGYWaepxbq
L4doWn7CACu+mpRjyO+ioSIF3Dud6neypHvHsrhrST43QnLD7zaL4l1Pu6/Xax8Tg421AOqg5Lag
PfHB11BJgOQCT5OpcVE500dlJNvIsOr6LUo65dwgAlGa8RqJFAReMFx0JPuzWJcoj2LER8nA1lki
Xb4QmCi/4rCbzCcxClCDQhP7vOXA0JS2QUPuf24oal2pjvxjag/d0oYzO7vos3PzklhHt9E9ES5Y
/bMQSb5xACPqGMj9HEYLYXeypkN8fDD0ac2JIMApfVbbd6I2A2kTA+eiXVzMIEBqt4IZGBgg/SQ+
6KiHUQYnC1dQ+bpE+Pf9CbeexPOGMSnLkaXJlCyj2akKeQxWntfd2P11NqiobDTjQlKL2bH0FS+V
AeTXFxS6oznFadGo9xn2kM+ki99MwA5IIdm+udKbtNlL65vsVUxv5RmJiPU3sZsJPlSlRllrljK8
wiIavkhAFA/trw7t6ri0c+RTpCJYXCq7/IGDD8Qzp5pD+Q0YUQRm/ljLKdKnzVTSc/gWoQWCMGXl
f0+wzNX9FMaP+nYalMGEcXaudtnCP+/WbMXMQVYLWFcNTKAdZkbBYAN+aAnAFvJywR9h1g0TL4xf
jqy8NU+/z35PwadYREdAeVX4Pk94sKz0kNrEtQ01v3dT2CmwhH80+kTtFB4mbG/P4V0+x9z2dDxC
GzNBDkCmHP2/7qf3xflCt5MxS2qrcxWpvGs78J+rNFQtyFywblhW5TEzJkV/fth6XC/6lLf0yB9D
n/I3Kkvwvwc+s9+74VJgVQESQcDVWXCH7tLR7xibGVWaoQBZKJykprWp4RDhgpHO1x9hZ86mzH9X
zWlme+6zXIto2lNieMICYQpoybOv76Kq4to0uSdRMxndDCCRJqzmhin9IJ5VhGvn3QSdJc8oRrFh
cru1J8Gk4rf0g8acIXNxWm4iv9YTJfMsh7p4akrz9SgUD7RmEOee+2rwj4FfENWbs7do5WzT0LFS
Jd1nozHZMX1ZAR7ShoWiyHh35FDjf53Z6igXltqOsaX6loTv69say9EW6k30Qp7mRnEhcKaKN1ON
OwYxhK8I8aTtBo5fA+ya81aF5fFWq8rsNHR+0SikBL5LObdCla3IafWsBidq7zaKXNz67fOp+T1R
wh6/e/kWORkkBzoeYXEj7AUhOXCIAulXd8ui2QV8Z0cE1P2YvgPY1VmKw8N991eqo+OGJgicMST3
ls+X+RmcM6RJ1pVGM7Kr0rlGfoiZhCgMR7VRdspzQpn4KpSdxCsuOgHRmxfZLIko8Ky2lS6Blm6b
Bvz5+ZiEdqkofOj6Tj5iF8MfAX8474Xo99+8tKia9J0IaNhTnus1LLclbqDuqrIfPM7vh4czrlpB
bjL0fuih/O06ZI6dUp4o2cypbJYZ6PXuZnAGqQgkw7IkRDKHdsrZYmgw26ojfc8CQAmLHTsAOCxR
57iSiaVGocoAFf1Spj/9biPbiPtITL6WmEfb3dGrpN0qX+ZCBbBSXqzZ9bp1aHagHwfVCsFMocuM
PyFG8PdWzsX9VDDjJfKIBIljl3gTcEt3/0nTjMukiRxW3aOG0dtkimwkHNmc7VZ74rOzjTwobFEd
7ajdRS7DCRmucW7JWpbfUMoepN6V3z+JGTCnNlLyLsNEYuCKNjvIgLepmwunbYjaUMX2cSrWGMzY
35trewXV2/W2k459+4VJ3Xa1oAwDsjjuVz7BZnJxMsqLr0wvSmxoOZRNIbL6qtDZL3MfenX4gULt
ijjaxTiDIz6iBycXGEXqbsLA8kgVia4j9Ga4WUy1YJNzFSV8v+UPKBmorXuS58DbqVbIFQLGZuwS
cR8aSEZBDODnLRgi9WcEdvmQ0j5WoSd/PFufTlFC0AFF0OgsNzy7x+S85sTm5Lih5+T8ag/wfDFK
CDGKzt0LJTgifQcsqb3fWP1m1qLq6n5H4Yu7w5yXeTSvQxxfO/bQy0cQb6RimYfDoQsfx1Zc1gKk
TbL9Np36XfO1oBSM4SuCR+6JxSOE0uunzo64ro2W+AEukW+NzVPqLVFfoPh31hCEv3YHIRFfmPCx
I6cRtLraBqQFKEXP7B1Fm54ql21lXHZgtRHyFysgCkEZLVxgDY98yPRfR8expPE1+Rf2MHDafQWF
5aj73XMPGwogpEWv6srkbKL0rLoBesn5mojD2A/aUTo4YA6ft4Y/g2rPBbmjIVFtSJXpiJyUopFe
+HFPv9mdMtsJuFxJ5m1c8gMcVcjiWFbxhUjiwhz+Pfxbjuetif6MDclsN9/dbmcUEQdp+lef0FOz
93k1jJB11Bf6zXlZ2x8eniewyg4n2o9X2qgCYFGQyiGkPvM8isMhM7Imd1xB1kXC+t51fQ/zCnf9
qzqP7fcfQXlEc0Z9XHU4f606qH7YSOwCh7ybU/LoRqdGsQQrNMhWOwcdp5AJxjTv4oYJbUE2LtVf
HE96Fi4wQPLH1gVnWYfD9RkSXl9sYtkIJCcB1J4VTx1Jw77K47sBPCWmQwC9gJ/ig1q8VKDkjhG6
HFs7YU3AoLjBtK/HJK/p6pgGYxuB3IxBmKO4FAodIwoAhQnnK2pUEQVmZTAn579CP5wDSgdVnonC
1d71sEyKrI3UZr25ddwfdKx4xYjsoprMYJTpTN5kHSb+tVsvLDiJ265DokVzEjsWfqI/sVUFY9U8
M9usUg77cTcYuj2/sappQinaVQ5yQ1PoLdAMAgCj1u7T4RKdHTR5hH204XhZFTSnoow7qDheKuXK
ZQVYbF4BMtEGRziZHc/M6k3pXxuLyZtmdpalQrrlnYCH2SKKUasGHMLVulhIB732f6W4WwW1EmzP
jVfSeU1yuqpQCBoITGi3cIeeG7NmC+vhoSqC0Zfxbtc42XPqtXgZs5W4wGHoWGTl3KgTUOkEXlpG
nYOJvpLxP3+EDrLPMpqoaVTPdijnlQT6WR5IX168/XBaXNe5sRoqyEV5IQyZyZ2hOKOkyoDul05p
5PoPz16zsdLMVY+l1OeoVEMbtF/MPyoi5416LoZcH3M7ZtVXkysovLTGyP6nAO8/XvGw5ME813Hv
XRI4smzAIJekyQixP26LHftwkZd48fhJ7Z54ME+qWqrKNOUzsHjTGEMgYySOCzWHp3W0q1/UU1Az
1A0JPB9zcerv2q18ElOcws/4QB71h6CTH/s5c7DJ+6hpwL95j24BeNASRUHFbUTlBlaofav3mquu
BeW85OCfdKBf40R8k4Y7gYqpHRtrosksLFXln1nTAcaL2LoUs+3opL9Ex/ymGGhp6T0/Rydvbz/j
x2btRmC3o7YhaR06KF9nYi/qF+i5ZSzWE0Mv45pcedxVBNPHv4AU8jRXygq5uhgya2rEMKQ6siQL
emISr0tHoirGbQWfFlp932Ry3S0e66oHyCwDj2wJCwHnvSe7i23dOenY/8c3yJkbIm7vvUg8wGp9
NfVeO1odRl8S0FP45zpJrDF8xmZUt8ltddKI7H2rfo9f+7b76bff8+4+GFFUaaiLcFj9pXuyYr3r
ufZmrwZACDE+g1mIjmpS9ZTbiFdGCfg8fMFwGrMX1QnYDUb9+F4ZFYOau343d4Un97ZScL7uezmZ
0hMfAyOnpU73iLeVaiezGHW2QNKTFCJ2JZfmrTdI1dvIBn0QMk/TYK8B1cMIpfQZYaMXvOS1idg/
ybq10T3hvsk8+Y/0yVBE2K4UHu4+4MR/5fg6duOv7/mCAukDHVpc8BMNjelXMTy8efTq8nN5WAjm
QeCiHFnD+19ca2k6rprIYZnI13DboDUkgTfsiVXI4v5s87svcbK6QC3ic26Yzg121D3x5yNssYYu
Bm5ZnxpGbkLGc0kGtPUDA9xHp+HVVhSAcARwQ9KuZ6lGIsTvLqAfvAoRmRXmnIWb1Jjgk9evqROz
Tmq0h1saYkLXHbvy+cgJKLBakCzeadBxA2mFQBQWHrjeOkqKTwvYaDrVt1gZFAQfyPKUpXfZbeFh
j/5lg5acL6uoTVNRvqaIrooCsKmeUhhYr4DdYin9B7HqL67vx+JHbTtZBFhKG/T3TyJPAH3nJU5B
8ITaRqlALXzswKqGwBvDPEeALIUeTW+vyzZRkh0a6PytDeqOwaO1tpscof2XjJG88LHeILymIQxF
fLhdjKMJKhon5xaMMShs8i0TLbvvLB1LsONADBlTVXaWOXsePQRJN3rZyURn9pP2gXIbFjQWMXBS
EL0+qiR7a2IGORQt2zG4WIWN5yVOZSD5TJo4d4DCbjhngYCRbDgpFlFwJn2dIT7VnXJt5l+9xKGy
QQs5f/mCpYnPZsMPF0WhLXeRGEfr2wfMbl+5p/Csyr8XDK+746i3Kw+heP0obM3Z3vlHagGIQN+k
DmFHCVepQXIa99cktAYydVKwbn7FKcvqaBuhkZY0L7Ob8WEGYyKib39YF0olanee4qMv6qCK2ZSQ
BUqTP9OTfG6bQlaWWLikrhHtcVl+i6dS2BEzTg3q7T1JsPDE1gzgqQitzWPYgFxk1V/bqFDiddLV
FN0WRwaR9fBCfxSLuF0Yin95NPFD/8jYXtT92zctVBSp/JFbefmEgZ9quG6XGFixIO+3hCvo8IpF
8K9oA1qvLxqkMNDHMdZkQkNfD6XYYn/XmQCMqZQgWCu/oihO+hhYxLzZmc3qX5sOYkuPs2ceFHEW
7WE5aVw8a7tVf/cDj0Uxz/OBf0H9cGIJPkdslCrKePJkoZGx2iS6/QnuGhO2UnpssOot5J636gsi
dD+4elzr09MCrw0BeJv1p5QSx9LzdNjY8D1zUp0UNm/IPKns5BSXHYg0xdlU/fxj0WNp2R6qnGIB
KkyitCBtECTV1n3xJftlGFBCheg30G7oPWyQ/OPEZP3Hvku0e26NaJSKOIWNnriZAJDptX31AF7U
5X1G8TG/xdzNF7rEOPuzEOinWzZJ3ZXiLUispW5CB9nhtus3kc50vZL1GaI3osJo6LW1qmeO2LJ3
KxALcN9K+y4HzTpsaGYSkAG0Rpm3Kgalp6MIJTTQ8T5hp03Lyx2/a7n2DElGdGXc3y0WCwpOH4vp
ZSeYnB1WDSz/cUyDH53mlYTb+zCyPO1UhNEqvWnCF+XlZuDuCUZNOoRGRS37HNzzTXB2cwE0NI6s
/YXaMN5vWRwjfpfTjRVr6J6B192oIq2YvWdoDz1ZhG52e8uztY3ocIbxQb2X3pL/xvhHhnDyfUsG
BoqCQK15DsMZolRd4ep4jkKenfkRmrAGhebXAf44FhXSkgRfnv7OpbzK7bYpmbCCVv4HKQEam/T2
a2LZnuxX7pkA3D2SAYfrZeJCm8MPOH2J8M/CJgBByqlpbjEU9eSW4jRm2HBPBeOsEMrLKDpfuUXH
065kMkj79E26fn3KOqGx+kWxbzgJvGm+7CyphI0c5L7ox6XOU834gP84h5SZPyK6AE/6RAfjS9fA
5EsKNrAoCjvcylruaiwFltctJH6T/wpzdX6yKZzuK1B2QP4lTO9cWVzO+UV2xYWpCQKAXORryZT9
ODIQxQgBp805BjSNmOZnNyERaLIz8g64Xq3IlaHJrzKqaYLKtA5rSfitYt0+WT2mwogkj3pwWFxR
pd+MWxGF+NdU9uAiiqOuG39QD7gGoPQ2W5mx7IZiCT9NLE02nRh1YuStA7YA1qAVV0guMzOURBBW
9aJ0DdHWFpd3ARHnqomM2VQ36SnjURPYimQkM8A9k+tRyl5zjEZlLS4CENKr6yrLmmjomrj2Z45h
9PBhQdARN9SeJyJxk+kwC54ukGsExC1YuZrrYsHAdwgZjvbezKFa2rTi73N08jBrxq7vu9WyNaFt
mLk9UWgIMd8P3wHju1NasUWaQA6tu3hYefZhW5BPlYWVM07y45JQngRJm7zkpjMpHeUV8vLEV/AC
Z3vmL+RFgld0x2hG8fEB3AKtFrEq0zm50QAo9zQdJSUbrHFUKO15ahXovz5N+BLrrecs8j7QlK04
xX/n4dmv7he1QB1TU83drbyc/qbf5gUVyzM4yh2UZA654vGRGIhBbDDFVLvAy4pA6SHFo6+qQbQ/
dP21LD0fwMuHzyLqd3aQNvd7s4f8m74bdDhRhB9A2mFePKLKMMyjsa6I+quSeMpp2ZB4Xeb1M6BC
IwHGbJP+SYL/uPcbzpEQ9f+Bq2oZa5HCUFYlTYTYLemJx0B+Y/sFe+A9PsjP/XNlKCt724xCtYG8
OGzbgG4qycBFE8VL7IqgRczEUozFT4gC1pE7VE1rxCG+yhXm501hkdrbQ3gxaqEG1O5sAnDlhNde
6y5O5+wQUXNJX7bEj1IXaj3E7YrmiGseg99wH5rGjim27UYimCcBTkYjxDQ11fqNz/c4MiavEv+e
CTBpq3pSKYndygzytasd1jAuCb1RFaxCnzxSwTBBLpWIr4rCOJ4a1Z/Vinf7VcnGxoVKGUHfsZt4
6+BjcfhM9HDcQoGPCPrZ9YRaSIl2v8jWc/s1/qdkV8Ji7cs4qP1E7HDyJ7s3IXTqGnlw3XRWN+gw
ZDwK2MOWlG0ThyJjvBHDErA/28y5b74tLFAN02i+2rEAzO4rz/GYKIYPTsE8Wt5mjWTL53MYosxB
9lPfmfM+EehixRB+NNrNbINI1o8gROdSP2I41zHOySANTNyLOgwhecybLPNhSGKwCZcW+nRy/rOq
/AUoCTXcU9oWzUcDcDZ2BHXaNVouXQ8MM6oM/6HbjGfLqdbn4at8P5gg7JDI6lF9XFfyJXdD4xQs
vMPiDrQ26as2ZaInfPOJ/lntw/Q1UvkxK+XEcCfninKFgXQ3Gp0zGmZaUWu7FdNiq8fCYA4tdhVZ
0LgvoM/694urspZT2/eA75M6UOgAkXCr7i4RcQVJHMrCpEKWHdf1MdTfTqLzkF56nz6m5iycwKKC
dIQ7Ff3vfefKaf/EcquWsHAoW7l4wC7iuY2a2VQxnFg/9AUxFyB4sI9EM+qBbzfSNfTWH4un5/Xe
UcsC/pJl3h9fNJteCJ2UXdR1Y9DwRqK8zyx/VRMeZTCJrLZ8dtv+BKtGwiMEaVdmPSuTiPQ9O/r7
6fuxmj04f2sMC7qsfmapjm4e3Ntj/C0QxP1S8IGmgPwC7ZuzbL/3N8YjH1WOYm/fHGOgQMSnujbz
XnGeoDsDMbw53NxBBTv0nVvWelgp88vsfs8rxUulBRpYzIPw+pputfpMYd1zjv6+TzbdjguJma48
Px8zb95eOtXFvStB8Gpzz5JTK4B4c7jqt9S5fTVSOkKQF/2BmJujBy/eudA7kL3XCYRTA8lRfIHO
3/z8YeU8ZJ3eRyWmMHwjG8bxYxDuxUe0IC0QMWZzqh2KVNpcYHXH/HzURb9kK7LEI2uSoKKhl4Fl
ka2hwJ2LB13Hkbt4IVJyudBNJzqXTfwlGahDtvYuXUgn4j7krSYy4l93D1I40jhOsG49eAnP/aHj
uScEggPXiM5ycpVDs1fWvaaSwgziz4pv7HQIdwbOoUzcCBO1GcHBg3ZTlTR5atcxdI44Sgf6G1dB
yDvAk8GCV9bg5nw6aCzTkqENpsGyndeeqPySPQoDXuRneCNjFAM+Xw1OpH3FUrWTkATeavVz6s7G
w+etsM5vPTWyQKfHzzPOSjBYchrpSUjGTj3j9oCoCePhju7poJK2txWTnBxNvJawDXIhQ07AMBlP
/bderH7JOf30JFVpHXzbrb7EsevzqQBHQ1HlyID908W8yMNSa3bGY+Eu7CXJ8hCyW8OujvwLA+Jb
2phw82e5AHnB6wS76F0QRzOCarrVCM7RWbU6JkTwJZlvn1OOtpDY6YXiYqKPthiRxV3pJEMilj8n
TMwP1NhGGB7O3LvMSTiqBt6LBwyWml4bfN/sG8pz/1rhfG7HaMG7nlrm0C8p4gAMxWMOhRkvA1Qv
jUibCySN4MwYmdvumSe0mKUOAducycnnZ5veP471stbK05GdJDEJXxg5uq+DmCtcX7en3QVGi93Z
zAQnlZ+B2WojnRdGuwSxy7mm2xMN0jrjPXVXk3W5PE/m/3DakNMU8ty3xX0bSS93a3HcGtkZOgLT
k33RG5fKM/RfNX7ZbvcweS1JQXIAj0Na5uwIB8XcIgm7tD/eNim67R9JZtU+aw4oDLKqHcarhsa9
n8gYNVIZGoqBwzpUUOI44FBJtxMnVZgsMgPu83D5hQY86LooigHztiwbPXFd7B5izwN/H5aMLGxO
IiJCfUneJQFrgB70lqJEbT4N3ekde2x99r1SMoGZ+zOTVEMk8vhJwv2NHIFSOqRUTE1ku2rItp6g
jm6+QmAgILmu0h/wh2PEfbOhDaHGofqVZ6wqBnBoD1zK4YzXC2FbU9em61hJQ/fbge+ZghIbpFQ1
vGxgIMQmur3KYCBk9F3JZnmreuCZdT72ZoVetbJg0gXKYf9P8KDYjFr9KSofti+c6PDA23VJSSwO
hyW4IL8xrA1a9O/LAHIFZcRfYIHJbO6g3UA5hyDNxZF9gcUPTXmQnktbG/uyaFyeQbsmx5Ux2Jxm
b99Wg8GDxb6nVZ/BvAYmil81HIrB7mxUhdgJAf6WY0h7idM1RBIkBMbvuMKe4bazVugGIKR2ZHac
npvdXdBWJq8f9O2MSvGFlcKNrD525SULPqVMPv3+2DnaF7xE+PeC7I6jb9dZ14si3aoznI277/1U
qyy2711lhTX6cZkVDIoI1QL1bPXZDSi1yWqTYAKjwrYhMpFrRI8Fxor6b4K06aQNRJXGuXx+mjT4
gqgpbTnQ80G8RMgRaUKxKH7H1+n4+cdmAGAPmlzIHHaGRsmyUSPL1TMJBgqe2yStgr6EGlzbKzuM
lDv8joy+TyTPDDpL6axJsZWo8VJn6LC9gobHI1hmyDfFT5ds7mJgFD5FQS3MPwrT9CGJauXabyYr
SJxsLZM575yQrsx4pQqBFoalz+vfM/KKHg8Jg7g+p2tpP1aBAipLAgP9aSPsq92i6sRnwR7WWMYF
e2zsjSoE4zklu+3ViOlAvGhxjqFWbFAEuf+SF5yUvW2Ddq3W5nviGS/XJxvAkwBK2iusgRNRIHK9
OTnswUeyGr3S+knj9MYBFYt7vBcU4pDHAyjO3sR35eQb0p3eV81gvjjW8mQJ5XsRN2zXqVWP3dmB
NHtFzKLQSY0hgZN6Co/2ZUG481mGnzrE9u5UTmLeavkXoAFTpbsbXTYm6uLCTWLYH4N0M0Hk5oNX
aOZqqmd7za8Dd9lYuRmA4af20R001TQACJIGvtkVkTQKQC1W6JTK997GAAlYIPL8CeJnLTyF6oL6
CHVQeLzaTgstgEPO17K0bI8/0lJNiQUMOWBegCCCGf8UglXBzChd6SK0uuJU1sS6j2WBY+UI2Q1M
G9xVqCxWcsUSaqgUVPpzEGVptEgOi0sNqQ0J5967QSAHdGR3KTlLWmyrMXN35MFhoGCBIERNwZAk
WPoOcHw2sr0+1CbPIvTfQ/S+p2mtx3vdgJQTpcfMKakiy+d1cxmgmviFrRNbsaaLXepka2IkpB+a
F9lkuzZ/2CQosz5VecRmCljq/zW2l8UsE47NhSKxcSYWlWTUnUaoRH3nfNH/+x9DF7KTbJIaO83X
5f2ZqADU/gQGIFBRUqA48OycAuJqvwsyl8SsjJ3qFiYHRwJhHoA4HavySKoklfRDVfEmrahxmECo
/nwV6cGn7P42/xY8Hgvlz30hddL9ncuRRTgVYXOu3R7cKuyd3hwVTGu+0KD9iLwKqS0YNpRyWuup
0KTf/qmUjyfPDkLqipETO9g55oj8cxTtedCIFbZ2aZrBnnpe+VbVPtjGPrFRLSakGdIyRvQmJZHk
aIv8pxJAIZ/q6PHNuiKk7ReY9JAu1xfktx3QiuwGWGh5CAkLPjNVE0tek7CdexACTm0TVUsdQeS+
DGQ+u50iGf6A6Wliwsbyt027PBUswKDK84FhgmSoX1aG1/yDr6/SWnaVjeZiZuSaBN2ijf0JSdSP
Jj/RV26RcxCc4f0EVyqxkVO5cETTasVwbUci8JfjMusCaTbTRm13WIkedUoRHNrbhDkZ6Bd+mpH2
RxROqt4SqZE+IP4V6QVwBuMl0xw6OgrP9GkiC+gSGYEU4xZZh1KeK3Qz2gnnYXnWgqs6Imsr4J6E
qAV6YvR9QA16B/E0E2U3RpvFK+yppjhVMAmY5MgrXAqb5OAxdqyuDHLgwH8ikFOhquosdV2nsDYY
ZqWLGdhAd7cd9Qt2uZFIKnhi3G/gbcuc6UGe1rOJaXJWOUIONtgjYrqdVI7YOJapKiI3/RmFDgSK
LWoaU7LtAVKbx3lcLmhTab0u8kHZWbK6nVBhLmGIHhJyfS5+0B1wRPOkPo53SZ6LL7QQega+00+V
xpL32xNhDC2sqflJCSWISlqgFutpPL5g2FJxhsmW+k0V2ske0umh/leK7Nu3hW3buFRlB4wVRVNt
gSe9o38LrIs9JyuRzqnYDDuBCjFkOIVe3CQOhFjhiRV57cdBThauhBW5UdtzCXJbEYzKU7c7wM46
4cGlhj4wDDNsc1NyxqrMGSX2vSuWgT9wW1blS/tG/1xtms2AY9ivemea6TBGGKEybujp3E9d6WaI
FYHv7NVqEXUHOgR4jRjD3mDEUx84jElXFnnSgC7C1j9MGgR5GVoWlY2/Idoq4VJwUp3L3I3JtfKB
/8gy94jGSLhiGzgQa0Tq0qV3NgwaeGl/zT7l2e2gHLue9HRA0e4uf8uqD6fChEm9E9zf/mpJ6gLv
ugH5seipi4xPNK21p0Fhe5dsO/UXIK8Ul4cy16vxYePscSxOvgIxRXEuP6SeJfUwrzaKxqswB2Sp
3JneM/KNx53S6nkVDb951mUTmnmG/JN+txkBMHksA+iB+37cKJuC0xCmLgLYkOEsEnLc6uAWtGqq
W4RrT9HxYiYAfhxW9Oa8f2Kj/G4D6ReL8w/aNNC8ZHgVsDLyU4NbOn4VDpz+bdVg4ToD5utTzU4p
Phj3aVcBIjMMD9eKVv9tBKSPqHId7/VlepGhW4i8Kq9gr4d+l8MjccRK6u6BI4o2HwJfRFdUEBlz
orZbkszdQz0LXziTvD2oGguZRgAL0u0cplbYF0GfidPiaQS5BmSx78Ds0oQ3xcDvNPfODAjsIAUu
nRfm9j6trwa0BHwz46SJXwE9EGkdJ03GbhY5usum8o/BdAmeZ029h30D7NhZHCmzlKD3DXkeYM17
VBEh1ZfZ5CWDersraO5kF8MSteUr+mB61F3ct8jinpLG+wBv62O4pVIsP3Wk494RzrujlRPAkcP+
ZOADrrBWIvpBImRF/bo/dafceWrYYlr7dhYaWlC1N+yzsPfBjOlyfEmrCkibpewLIKh5eKWTboHE
6+GF3NjL4EUxS38zQu43/0zeW2xW9AosTHUsQnCPeTmM7p3122hBf3qzEP+LJwyjRCxWLilph/fa
VaEbn9c5750pKIrkZTp9QiMlB4R6Vdrd2EItPC+TD5JEbFQDQ+ErsrYi6XgdnkCoCLdwXA/nxonz
qiSXPVhqF7chhUDk0W7elwzi7USsvBQS6WDyKTpI/p8sw8XjLFDdotwWjJ0t9TTXze4K0amcJeG9
Jf4mH7rMkuqH0LeFWvyV1DqeKRm56zJ9IbBgA/dPqwi9s6JiJTI/6FXze8ltgMpfAJzf1SfQSuVF
kQqbTkPCyJkXy/cNE9AUNd0aRQHLfJsOhi6t6jtoPldLhNGoyVmNzqzHpRTFcAGxNkwerXsUF9F0
T6nWPOotccm0pc7VgqEJmuN2i802bhWFWRui2Xd4Sm47LhKunr2L99FM+S/tpDIHaSQG7i59QAVZ
Tigmq9hb08EDoG89Ag9jpZ8yBPtUH3pkuDt07AFiUrnCGiz7ubs0wrlKj9xPm3OEI+mVwEJWaC0W
sooTv0BZLCKAJj4IU6VgNJh9dkjfohY5p0qH9BGMDkt9dAjDZPaknNpPvT31u+Djx7mlFjLbMqIV
uqhIsGxXjziRAUwnbIG8Fgg2TeaFvQkiGUSPuI52WePc194w0P18JDRVT3EQDKHwjuxBYemEaq5M
g+6VA6XxUC0nBAYDxCeHG88Mb4dnJ7O8aS2iIPYzXSNyM5tDD1gK0nnh8CrkK+v2q4LBK88o5XwQ
lYEvwehTeJJzJjYluyPNqpI8hPOcaDLAd/29Ze/BhrAp3+Gjb+T9VgX77KtQCkWfr596Fhld3EhV
kgiJdAtxabFsJuNApaW+aFXYNNcQw5b7M+4yk7DqynaCK9L6ijXp35KOEIX9LtYATL6ZlMg5BP+g
FUjaInMIxHtucE7f2cUJ16+SxsmjUDLUNsPjGYAEpW31cq9nVwNIDn0cYROaffTKfxWRtDNwe79t
3UNztJBP9dSd38ZDOAsA1MtbVEcCEzgKVYGfjnDYAVpjTnwx0I2OA6enNkXSWk7f3uWYWgOYxOqO
jEplBHD0COwvGmOWmvzXeYZL4AkchjCr/UI+SQyh8nvbaxux+/41pKzFK86+ep8iCYt1DlnI8gLO
retiCabv1iNSMkKujjrfOI7Lk+Cxjm7QxZ9lmKdGpKw6J6C7pQDHJd62YJ2eKa7UElrdKvMxu7ip
fBPEuf4wYutOYsuyM6XZQ6PXOKA9uVVxdeETTivSb7uDVZqZJ20J5SG/icGbl93NIg2fmIYoVTd7
Ckj0ifs8HGC/TMlzEkLh52W3ed1YFs0YXQk7Kf8n7uHeg8LL7LQ9TUCr5Ml/ueG/7nObVWdO7wkC
IyJHiG6V09KJNFd80oe6iz6tk0Ex78OX08zcqQsviDicclhRl+VquEEZB393D2zqvRozHuaGC9g2
3TuvxRWwWd3O7ls8Of6udr8jD3+Sf6fHcJ8tE/cs6WTRVDhXxpeHV7Grow7KTek4Lx577eQ5fTyH
rFLgn51+na3/ilcLOXr4JIyLlMAS0fdpCVDVGo00H0CH5lnk8DQCxWM88PV2ugWnYyCPRlU2UyXR
spISl0Ts6jNkEEKxt9i3GzMQg/8ukUDeYRAvWXBtcCab75CPe5USr9quvLRHafAbD8OeiEYjBmqa
xniCs0zocx1H3mPZEWCMijYwISkBCh3dBEPX7IBfH1CpEoBThw1O20o5kgKZrIRmyT9nSclXA6e5
hEv2GFcOIgWRHNcOofRk3iKVp8/id7oBwZa/iyGtvRr/tzdQWT2eLf4xZ7ebhxqyW9wC49tuYF9F
NDu6idF5AAPAco01ERgqNcqCNU2hAPrMBPpN/efefK3WBXUTELZc0G16UYBID8fGcbwwgrOvE2t6
mWWH1p0L0RJRVWBOaCdSO0J+xqyT80viNMtsLrImWphQZPLOGsPDrTbcBg5qoVTL3ZpAQ+Pv7bh8
S0INZYIO8kVYA5HylbhijWYZ9l+XyhUt7vvhNe7/QGoJ7newwapMvC8cssIe+3V8KN4UIFLALDyM
9Lhe0OtiNj23o0Rp1MafkpNDzLtcWP1AEvH2VsNZAd92OPSAxpHZ5cOaGFOTEutIlOhuDq89ZqAV
eIwhoVALFLQN4/Qi/aPusaEivKtr4SI9F8dNZeDJCCnQBDM28ScsIUKZrprHCB1ikxYZrA6+CYwB
srbzONNbrYVEms0K0bM2FndqGM1gjy3ZCjMnehy71CWXkQ2Wmi688GMolGwhybdxurBDbXqXIb+N
Vm7yOE9Mm9aVqinsSXWTNpun5bcMPHePDjUg/3mnfqhSlxH/AXmIDYWTH3259FinyH5UG305iplO
b4tldjonAuQ9P3FcKgny69OcZlqwE11y2dnKDkv7runuCDW5eb/ZQ662YaU73Uw8E3wQXa302PUL
2+OgIDKbXdNWZ/lRmuId03mYRUa5GDJozAgQwhb29yWnrDCtteDvMJdl/A/nOARq1FH7qseLQ9Z7
ss3jN5jSMZv4upFPERmd3idT4rcSNkwvzEkTTQGk/aZCvYeCWmjBitIYKhZ2pPJ6LBIm1qv/VFwm
qfBAPVLbsfpUOscx2Y1f1yRtnrh35FAtdwODF+a4VZU5XCx9WeWyb32kV5btDL8cL/rKTqgPMoEO
vOHSKoD+AeWEOFLWmL5paD9KewX+h2QUhwEoN5kMUAtleNYXje532tILutrIcVnwr3kdQMd3XLqs
lDqZb9Ra0730MYwwwaZ/5vGa/C4WokAOs4RDCg1bESIjxl01cnIIIPwH4eFjFPFacVabI9kBox+C
uNNlzcNu9uoPX6qn12C6+tBpqrYKPTc7YfjwmNx2w+r1sBsIzd4yU5SEP/80pZ5u+xsAGOCxX9qr
pbKiTgA45MptzK4Wh32i7gIQ9a8N6VQQDu2ukH1NYY6M2r2hzRlZBo83X7Dwr+0Miu7DOX8izoSV
wWlv0AgwZKJcYNcXD964q/uot07d5m85Sg7ozkA19hMwK2b8Dxq06Gqr5uv3U1oU7YM3GO7HAFSe
hsFDORNDIusE3TP7Lx+72IPjEekGy7yi/BoWRI/HeRVEWGJQbYxlLydVla2VCpru0EUNbxl651f4
mwDM9hFQKv0Np8GCWTlwr33jK5m4mdvxTkX25is8m9rDeEQ+t51cUZUME63pOK9NFBya65dxP/tW
/TYXBxtAWmbp1vhPVxerSMIOzGJ//dAH3YnT9PFkFL0KYzibqr8gOCDo7Xk0L4b2zYqxVUu7EOXl
r/wdWBX7A1tG6dCHajEyft//7IdhH5+DekRFi+0zbdj34SXew6KTwavVgz9HMZ7wafwqbk0fIRpT
Yh9Y3ieJXrlaRN4UzKyBBa5vsIsopEntw1uO3ZZ3nHHrgstWTjdEL2Y2puK9i6JC9Jd52rvGHssi
4ePJLiQcPdsew3+guplO1hCnceLDLrcTwshp5e7hrp9eimKwlvYtYET2/xpuRraKHnMdqaf+7wox
fG+4zRa19Xw+BLuzy4S5fTSfN2AUPsfJlpdrkqwAKM46e8J+/plZEPBwzveF8aojmZk+MccK+Zxk
AKoPaJsRQRRB0Oy1dNoAWQDMcYA3Jk7wXFQqi7lVmeIp+EGcQgEW/cFKN2g0lwJr2jBFKn0JsqWy
DxXp77Wvgbe1/NxxTOQyQGT6sVFNWylpfXoxngquNdOB0qfXLL/+XWhk6aRwkc/YkrU4E/UwiJZf
R8Ci9bxPlQIT86o4+EkSiRPq0v2vu9mfczJtON5mJHc73KRd5nIKf6Fq0ywlCHrRE5FHcxhcssTc
pHBMPs6SI1OMr+biIMIrmAnaZ3hshxfNTSjDxNbMpBWGlDK60bXUF3sDL4GYaLNbYz+5RgZy18bl
ywm5ZnUVf9yRBY/AX4TUlk9R4oOyq/+We+PZ81DowDjueexCpOdLVr5TDS+iEDxa9cTvR/1yBl1j
ZXB00huCLBXRzlbWe7sbL25vvxVfVLorXUtQzThRFLdqPwS2bFNqnnitgterj59hPAxyH6Nu22fs
zF6lUQDxcunmfsQP8XRmVXdpiGWQRxYczQFkwFIip8NrTeXFQb1IB0rg1X1y9JrWWSLwVfmDd+b2
EPe/RZxUaXXXPRFCbriK/uSSN9AX2EVSSoqLeSSt/C2/qEguX6HuKWMNCRHBWu8IQU4rfQARFx1O
AvtUJcM6wYfOWKK299JU/Z8aMDHduF4nlBmMNDWNaiw+tL7aTbleEOZJGX6e72EJ2lYWXEdvc5Mn
a4NHmfFFC8MHpkHhZn60J6rKCqBTCpHk1pZ0MEDY2wFJrBaER4pfesvRvzPtA3SXzuRuxyukFbKW
xP+YdOR0uEPn/GseVV+oeRmPRA6N3Py46G7WxKVnztVhBV9sy38cjjoQ3uVo6UaiAA6BwRMtGxnG
ejdMJ3nzgbTF+fFAArwEWhm83jCTSo6gEkwwwU468hQNds7l0N6XTM4vGzxDWfs+zuBukIK7Lxjt
9ZZENL2I/zGMI/cU65G0UEMYSYbFagTLRQfuHW7K8pYbllD9LxR3VL5xu9B15+iIr2/vM70CWtHG
lmPF1lci9jLdgyk+lYNPjn2XL5T3r//dqzX7UWXPmScpTxhxzRc+2OE5THje1xcmp09Rq6kjceQX
kFktfz4oauv7bPyh2iWcraEZfvW0fI8hxp5Rrq3D2zmxfVOF1IjW4DzFIDVC71JCJx2lDPtpw/QO
nlO0L8/+gX0DJF6z5wAbmST+btyVv9DVOIRc79KYXkI1ZzeMWofv4/ui7xmjBowv5o+5VRkACRVP
6iAcSFq3wc4E2ZqYk0gu7xqunxxt/3NWTJk3PT37a3Wm++g7JkC5MJHf8SSHoaw7QNl7MZfbt9xm
aQlzwaXaQ4aPx9IKXb7pbMfBUZeRVr0YzXEjWlAoETftIR0dePVAGTogd82li7MIjA+vZuG2MvWX
lLth902rq7a2qp69ugNQdQ6VPSInh8whxPd2x6L3yHIQ54wS/csWClHVm/ko9K04L92rIqmjgfDj
b4FtHel6y6bT0p2pT4H90glh4jqVkaHKwGaafsULMWxgswp+yKomfgXLQpVnyK4ncLvr2gnpmB9x
5y4v8G1YUa5X2+6pj8nO0y9VUC/RxwlstIgezu+MhANotqNUuQUtULkJGLgMIXqKf+XfhSNbJCmh
clypJv1JFKXJk8sD7jPfApioXS9iU8y6mR/GdkJxFUhWLUo9TeMslg7Z+Cchu/3l+Jp8scNjYNUR
ImpP1fEI5q6NZ9sFBzehMQ9D6z38wgzH1Xo8LBBRPiL5X9tv8i0dbKTKQ9Fpu49K0Y0RsPp68m27
mzMF2Jln7b5XY7itiR4ZFHJkOrYRUIEbbt4oNyV9MMWneVR06FD8cn5r7QyHPXmfd2FgYhOZBGR+
w8Hr1AXciB4rxEYVIIPKPA2eARatH9T4udnfxAoTEPjXHjybFU6920Y8lN6r2/uMJS5vK96u6ucm
5fo4sOfOFFtmpqx/BXMOYBTULNwNT859+2woQzszAtcNJsXaoLxJEp0U6jT0jkEaAcQaBkkV+nX6
x/6ECNo7sQhHHAc3j7uZMHpsGqCk8TkInDKe5bt8Tcy+brRlzVpSy1AypfDPGXsaKRFcRrzDWGcu
4DT0sjXfandMfXy2Og+TWt5VyHVn+oYsW0bVvdKcB6LgsbZws+B75QBcFkya3wbcvCVQHre7QqDW
iCE+VFqZXpUNH10RRWSROHfj7G7/5jfH3qfLWru1eoQKFdADqV6tsuwOyI/tnX1quPrLMTtqof7K
VWeEoXfgMNZ/2Y1MFsLBh+orIeJzPAgLHwnh2z7OLp+kHzmwdxXaSZXfdIA0QarLZM4WqWdMUw6L
FOz1WEFhOVu2C5Gy7HqAU4X935cEzRDQ82lTEU8JbI3xkeF9e/BsZ6od71BKclvGbkimSVOFu7fx
HvEqV9m/UxOxJDj49vLbKPlGE8sH+d66xpL/mGrG+Tkr+ETtMjzuZgllFg3oyqBytR9odmQAP1jJ
rfzFIQXjaGxSSWliFV7gf3EpmNdr3EFN3mPCzFx5ozbLLtFHKhWnKQV/yHGqWIV+Gs8s/E7Y5PGZ
sJho+oNt41ZWCyeVF8xvZztEqR/UguDnGoF63JRBOJUnvhNDBjSN6ttzaom9hnOg0hl0wB8h593m
i0XzJ6lEvFyOSYJC5Sxg5b7prkAKugfTyrbLMMiT0rz7n4pS2zO3RXIEGyzegZFG0MJxwmCFPvSy
zkI2TLabtf0TOYF2E82G86MaB7Jkce3QRmAvme6MqX7r9tH7ZLrlGJh2fWTMZNScBvTmWDSLukhL
FmQgrxCKk/2tOGtFfzpgEfj+2ceg5Vi9hPoWdTaZJeYw+QYaBA0id+Lv/7gbawyuDF1EpQszetC4
iS07XwrpPnQK3GnzPrps0aKtG2ysmCu886bjwDHcGBrCFkWd2FSHiKAXcL0OAXUbAaSd9zJipbVm
aW6G5mdN/wSDaYaqtHXC5voyWwiql5tXXTtiaG3GeFFn7X/NNyI2EzMc3UNBNf8qDDTbPbstTb/B
0XJ6LXDQH/zsRXWDlIsRr0pz/nvJYcl5Vt2H3HCb5ycsNh9waOql4QDaZzIczys4muDS0n7RQRND
dpYvBSFPXPnZUiah9Omg77y3wQveGPVcAqWBRFOelgdYXwBAAydB9bMagDYLP6RdBqPoyJ4pIj74
OzwemCxd2dMDpvOLaxq572dHtOGURs1FpYA6fZYeBJNte0oHl0CMEKQsVuDEglHOYj8/Jc+fxdkb
ZkTrkI98Qoialy4gRpLJWtNpho/+rXasuXk0GWZGUXTWaGLOOBAzq/x/eNSHNxGUBFeYBD39gA7f
F+ia8IfAkg3zWw8FGHb0nguLFPVzpSKSa3pqmSK2iN+x5Spz35Ire4L9S38MLTxZRCnDAwkP+PnY
vpwzR88+RrIEc8BxVpto6A9FNZehcWEs+myan9BoJN+lUFOcen+4nyUTDgb/TDDdqcvVWT0XJjLz
lNoTICpVzYPio3MHsRLCP7ly5NHHcN9rkH7Trk/6HemO5suTOgKOvJklrSmP1B+K9OmFGy9xR1SG
SgpWFO61GVx3z8U2vOpH0eY1yLZ2zzvxS1l956HWR5nSzYgurtl15ydu207JczeKzc4oq5ALVmHS
/sGHfXwP3oEHYsCfTIawPKkjBY8/YqqwPbCGyrwt+8j/g0rW13kIUmxFzCUEaymSlueVt+ErVhZN
QQJtea8Qo4h+Fnu1iubAFL5pQwB3e/yjI5tIHRicatemcTd58eLocmqJzQryDzQpyLtsvEvQCqxL
Rsav+XHadPHnckV/bTbx7PzRf55Q5zqOe60uCLGcahhlPByVw3ZHJiHaRwElQCKhjtS9jxAl4HmB
OSuGPHocrT3IYquv4zF2FhArX1TuX0qkJLE+X6QGZ1FQgfU6/SrbvHQShsoTra/3nF9oqg+YdxOQ
fiDH2Fmgh2ltFGf9cVirZ8wb5VUztcWEbUET5hFT27/gjAgZTaHewSyRHu6RazIiW5c0qHmSkMVE
y9BHRi/CQ2iYvdoLIUbbxeLt+7uJoo4hvZcZ/tUY4YY/lb4ZX4rAQoj7F5EO61hJjnYqmyeRyzrB
mQQkJo8ISQyWYGNFkO1nSAdoGuj5/nLJjbAu1LoeojSIosh1vEYdTV7G2M6mg35Fotkv99c7c7mI
PuPT6FW3iMvXaAez+ZAJ4Z4yMWNazlWERoMVaGEqkXUjN3gGzKHmbUBjfy90IcjAnozp/lo7vm/W
gUMkA2XusyKvUb76m/uTWuSR3/S2HrtBuwoOIDfdc59bXJi8bjeUOZnUNn4Rw9k6Bc4DbU+FECVA
KYCI/RIdsUHaw59keCpdbqu/GMmwGRYMn5tSvHtv8iYneXV8ePJY0LrjoTrOns9hz0LZfbpvia8H
pqZ66aJWoiJDz8lIn8oLU27WywXuGhllA3CoBu8zD1HZ9zhtEabC7TnbVXKc63bLL6rk1yomhCi0
I69gUFmJLLyciyfbY6Q7oPrxM+Ahacqr9Zvksgnok7cHUx4hAXn7UkGtKtKRRETK1LZqUDVwXu5D
iga1BxAmonh6dLR8cjZ+i2CY/oiaksflqpP5u5RCc6mvngj6uL1HX/isot8zlinDLfv+JCP/dC2v
Zx8eQWV3ETJ05DjaTlwXOQFsvEsHJ4yWbPE5wVA2P3899iUnR4B/z8adjKzlEJAwKkXxURrAgXKP
Bnvv+z0Jlhzrn0+fjjaxAMme6hNoG54XqGhZed7i/77Gl7gUzdyIdEXJJrM2uPXqEJiULJRjRbOq
xBKHPmE1WqjGNbhK4SI4HCYervxajM7znuII7GQOCxEg17WpYMozUhJbis8AcvqX/xBrwX90UwiX
ycINHDfPBsATjy5WV+IAsml6l+/uj+gl/auXO2rbZ77rDqRXU5Z6dmTj9ZsLf1LtSItikzUAQj62
3n8oJH5dlyq5qzOudAyxwQj5VAiGuaKfAjhItkN4frx98otH0vmb6G2nHfnDbZd6C3+1CCB0HjNK
vPXLUwCPeC1lctvmNpU1DoJmlP+yb4MHqORejIlH7ZYEiwgzmhYGFSh41yCRcGzjXPL0dq7ctIvx
fQSEomzEwSrYdc8oHIUApWIucCw/45e//hxrDN1tyMTPKrPTB0OpsLkA4Igv7lE0JXsc3dk+XEhb
uPwsTophiDZpsQ7TfL7biByrO+tLq5i+ip1UGwqzD363R4HY8zWosWXYvikWSKw4c9sKlUufRMG+
tADOvdvE4q2xkYg51Ppw0OvecHEBWi+FfGwDwAwDJnwG87GXVt/IJBa9nAJ3iRYEm9ysiIAp8o9/
m2yzvN9XcWHpSaBNHbEJXetQgGIrftB7+H3lnXrckOA4zeRIzmH9FtLG4QJphsxux/VIGZwuXVBt
RJsyasQI3KnS0I7Hy4BPI7sKz/o+tShjm7upscMyGfQiPW/1BVddFYLkeCNvxPA+s+z5LNuQTyOt
HVMDGPUOsitgSHzwX8bGHpdKrxny/TW8mjbR9TU3O8+DPDlhdJXU+hUj/2mSRHw4GLMkxTDQL4pn
k9Cdd2O5JXE6Iz6CheIP6WgFU4TTl39AW2nJkFXbC53OV2OEn+gOqFb0KHIvr1ZjA1JrCxmDy3my
vMuCB0r98uZOURTpN+9NnSEGfhHCC+c5HxCpkTbfbkoiGlXccSHbznV/URX2PSLuINZy6Nr0tXcZ
esFg3QgaC/7FKbm722ioj0mSVhcnFXZ4DeCkE9PLsLCOMRywFzF7S7pzVMwuUa66S1zC6i3hG1tG
N23keGWT78lCowJljQYyk+cZ+Blg4/mW/HVt/kxUGDFn/yTIYXs+dijnFLXyXxMYvuA9vFxT/dfn
fxlJZZFd6TmnkANxpaAesw7LbzUowTAKpbBOEugpdx7RvotEPRdNszrXQ15/eIB11A9lgpkwamcJ
hqReHBS8ZY4CYfpkoXAX3mr/HtkqDfR0minTxrMzGb1bZr6GP1FfPlQhlQ4OPLjjIUK0OtRrz62f
IReJzyHm/7dnUvAGVBOGT5Tq4Bm5oU/cNK0ETir4oDRN9rSXVzdXpmef9VCFA5kzBiVmkXxdGx5L
NLr60VvR/931wI+YJK7W7nYtX1cTTASOHsckc1K0B/FmFLcSo0SFZj9ZOdgAHUMuk5LcjWhzimsK
UA/l7ilGlsg9TGhEc11vf9pVG5jfK7Y+WE7UqMsAHPVGzRY5x+cbY1Fc8olpCiW25QJ22Xlwxw6r
VpDAsTzzPHN+RGV5cpXtwF+gUZWcDoK5Dh6qQ9d4icyu9o9I5YavwWEUzn5KgxnV1Kac+XrTqZfn
beCzyyGkLcy3yHPZ288HuRVq8cMzbgcAHnNWVTuErh8nzPsKAacjFDYS1HYOAf6GZgOXWTMEMNGF
dyeYcEiR7DiohNPIZP18SYuRWhcqzY4NQGiLSfLa9f3kjLnZjESEYUWhNQfFlQguoaoqKcLhK/nU
An7uxipB5EZ1W7vd+fn4Rr56N2ACjZPVk4d3IFIV0W7eLvvMBi8FWSwGIli9zLiR6FZin7j0kQZh
7jpeY13c60Y4ANH0PeahyJ/hXqPTVubnnbY4kO0kIW4jQA+XD7pT7cgkwna49C4AQZ4+00LdrNpk
R0ShMaSrF0AjVlticsMbquDjF6JlVwptBABDxFiHTKuRuIkv+10ZIvc3SP36wQOo7MXb/0cI7R+f
S8r+CmcdwtdqdlZXEe3VyYRf4CYn8N68J5q+ruRFI2NyCmL1DOgdBLU6mI6pgZOqwKn1hoDkw6eF
Xw0VRtlhEU0XX6CtZMNSs7ktYFnXM7baPEpSs3+/rY4AZwv2IoFcuqLZWGcYCR9HVavYOYFEO3Rd
HCNV6wp7LGKS+JUCaONznhMXYq1RvdOfa0xxU1e1I2eH9gjnyjJbHFIYj1E2cvM9ms12M60TZ05b
jxk1SUf6PEEo0eAr1APT7oBROoG1fEPXVm6QOJkn4+zmBLnVvtHnVV3vns7H96Bp0cKIFMfie/dR
po5nHlPfUkJNHXXZVPzkZwNIe01EeHz9CobIOSJwCX5dpQ+F1uhyF2YXFR0ppAF4f7pRTFuA6Ogq
3bicjiQ169U/aGjVBpjbYovvinDfh7QvgNCMlLgj64xU8MGSWurPD2n2XpYYu5zXZ+bjBWbToUZP
gRxDZOivbYOr/2gUclca42dfVrWXqgNmSmr8pKFv1RYwqsk/Wx3IgztqByhnTXC6o3+Q1eC1ghEG
pYIKmYESoKQv01KU2B41fLO77EHwkmz/cORzVOfPIpQlknTij36i+xI1BF0w0WwDWzCgNDfBgUmf
1VRe2adnvyz4bzlRrd+kEmJcvuhtraVzcQGNVUavSwqud15D0Ej3yD8bTKW14yF1126ig2Hrl6pN
V+rFd9E8HAT7glvI10boWTa1HMEiE2PfHBKxI7M1oshPZwoaB/AwEO7h3XCDWf1tsO3XfZpJUi2p
bIQweAPD7caqTy1qmpVwzYWGA+36QnEor3veaUb9SJ8KwIVYhNWou3YCdUQoYCmTpBjwWoCKRZzM
fr8hrcScvmTjlbzazZ+nUptSlHokMVnaiVflh0f2pd+f0ojIHkW62OD1TJTKBoA0BHLiNgTsqCuz
drQwMIRu1sDvc2hfgqP+08xnhSyjw8uVMw3iVlvnwwiZlXHbyw3lYRSqgcpAOP28Em/rSKvGu353
ZhL5NqU0kV6BuK99l73YMtuPNRHGZOy3tgv9ezb942JZX8VtZIn7/AFUh5vZuWWpJuUkOpFUdX/j
e3LdbkqcCJrAU2cT8HRoPcgM+Q38UHY3+6AZgghMT6EP1rOoCug1OmYju/J4hVRiKsLDiJPuO0dw
cRDzbuD/PT6xNpEFaGZv5eask/8vfRHKCeFzYlRjUHDO40L9TSvEZoE45TePy06gbCiBXJfDxbjy
w2ikWmbmTGswwxZa583gjuahmNHUreoxftHsnFBIlZMnvV7qq4oK2xJByh1FcabQiEZxLxWWFCer
PuwHo9G3UUNtak1txfHjVAXwqRPmm4P+WgaF7E182NpoaTEZqWPj1ST/V9QnocH5uYwesZVMsx/K
P8mA3tLUhgj5kmwT9TDNCEcYsMplQLJ4o/B3C4haGdXxlBjIgROcUWOjIT6tEizy+hOkCLnXkjd2
SbuXdUIB1Ox/NPSLHEdXiRG1pHURHqvt4vanlTTcrbJLF1EwvDtLH/Zc9EgJh2T5E9a5K+t+pY+U
5JN11tIl4SpMwqEJlY02dssFctoCzg6+eFy7s15brKclSnr7SE4ok6HUStBUnNrHwnB43lu4iKQt
XzkWUY/IIiFqesuwtpEfwdj13OEz3h5QGah4O5+242pJMFzbzBI4IeRruil8BGsPd+5WHeWCBvbX
8E2RqOceyHwjy2FBTbMig8K+c0oxwNuls8HvlkQrT8o+4K4dkPa9m97ps5oC96Ql029s5W//9v5k
kI/WrEvcQTtj2jV+iNrturt3DvQShyoG5DSsfeQ0rFDtPAldzMNrgWdKrpu8v9QRhMEGW0XAOMpj
kgyBDKlERs4HW8srx7KKDM4CpmKEQkCeYfPrH9R8KOO9OYBLG4mrhKhi051xs5khQuXA3CZY260j
qjPmf/lHMfeiNa2Eb/TWhifVGDuEEdUpAqXTW9D2pJl0yp0gCh47mVEZ9AOcEeFI0zamG5mJ3B7f
8dgL2/93StqktqBh/66RE3yFXq2AmHf2Q1BL81UTqzRgorXRb0UUf1Ob+w1miKZBRFKDFaSVHEnJ
gVGVR5jaJPP+o5IXSmJIWhcqGq+t0uOEsUewl1e0fuC31TIDzJ7KhOymVh6VJosCAc7FH7I4zz4h
KSXd+FJBPfSq0vrfdPq8KnRCoxeHpH0L8NWTfvVOsawQPNXcYwLEVCcMmIRYalSq33MBUwfcXedN
Ygv/g90IClscbfgtz8QG8etiR+HLTenNjhHYTeJ6FP3lYfktc4OvfveehDgu4A64CrITP7Fc6Z8L
ZqGw1rZitAwF77yy9PPp7qnWYiyBvuLbDFcnSw9ftxSUZkHPyXFCr8cosAhLrsXi8VVzUH5qM3Wj
SeQ1KeDIHUD8wXsAAkEXpE2QIPPCmTfBz5ejC3Rn0bj/KA7/SbsZYOLn/lgmA4Ej3SJZd6DKIZoq
g/LsexzZmlP0oj2OEXoefapoyduj/EgKuMSClaxyv2O+u+J1D0CwNIWyghHJx9QznbwJpKeNR9m5
6qvY+R5KpO8fONMw+Feaey4NK3/dV6ZA+DyUNGU9Eidfj1te/pVkXcgawXQ+sZ01suf1LHY93zKU
akhnaVWAA8x865YMxkxdAC05CfjUkkxtBlYqjkVjCOOzpVk0e9+oQlljo6AMay5SEvDOy9XZOyvK
pc8xQsB2lKs022T9vSr7luJ3zQZVCdUBAEQ8CkTIVKyh/g9cBW8PJDFDsYq+srPED0Ez3CmrkIF3
PMT6HUkrJW7BP3vuzY9lFaqFJQINrLOrfA9fBTZu7U97OToLVK9Mm4q3g+93HL1I3wgA742u4vRX
N9Cygygjq8boj6C8h2NarGTes2Tn7ytxP1hZxzzKFM9VtvQYhchouBo0/Quw5PAHsys08x7Fcasq
n0k4yLVaeGdwxxkPTBGVb9K8v5tyBWOBxuojQcvjqntVe/kBRbnA9pRTlrdqaSVb3GFAp2p8BSjk
waEd+ELuC+ZSps7DiBpGtGw9BRefRqwNT7khylEq1bVUVyS51RzuXwSJHyiizoyYPkoNZO4uZZHt
2wxmodKIM1X3dOG3T32XWm856J9f2NNBSUHcj5N13mDZBfeHii3G6YAbVtnrtf5wmLJ0cGYrbvt2
wEs4k/eqY79atZuc30G95UO3xMF1+PtzFDttS5PUeZsW8FIMzyleN/UYHzI+QcF+1aP76uHXMvj5
Ju+dMIlB5RdbyBdRlWEjtmHVEt9Y5JNgwL3HNpwp4+8XcKW/JFM8i+NM0rllB1Wv969N28s0qop8
PwhoIXEh3pqEL6Y05WrK3R2x7H5zxe0m1jkapoNRWElxcQ0LDJSBcsFauN0jbi48APu0PzioEDNb
ueud2smn9PKJ7TwTkkoAM6Uv7mD7SXlux983Wuf2p05dZxBXuiQtLa6NffqdglJdLEthrrL+k7Fq
GIwh5JkoItAxQXzXh4LxCKPA5PkPJ9gL6KAHjIynTMbxmAiLEexNHkX6wH7mAR7DYS508aEJr+PH
mbF2vbGAxFhx8KF0K9oU4N0Ldjd3hAurqRULdceyqI4SnmoJywE+WPD2PqFAEQbu59U/Hr9wGHZ6
BZGc23NP82Q8RQNJIxJ+MPGT+ASHtaX+Cnvrxr5YltVCfOt+KLw92Ar4VsxCxjS58mlCHGjolGg8
9vGs+71NZeSLXgQVHNMD11R3ouB9JvHHjW8dT0hCAnbe6LlfJl9j3/XZpHWuu/6p4I+/iM1cAtTn
pbkeqJsVvpjeAlp3I6CWc6h8e6gbnDXNUnYNi++4Oupx7RtSeqG3KyKY0wm7/ddulOz4IYj3gFyM
ThjfrAmmqZmmGrsxxVANJx0oWRaTQBc+kq9dXTVWOW4o1gXGNGnwJDl11VxVpayEehAVvUOpb604
25Bp9rNC1pjKvdYsdA2LVKmDnRYCHH+Y2MFCC2k6AV/QOUXFkXikSTjXtKboXjKDHrurpcAJ1tHf
HbcZKOHGKxIFAepZb8gDyIP21VEMgTy24oehKcLqUMVe1MTVLsI60YOUSYiAhadn/BLmVU/P3xXa
WQzpkJBeMlGZkx5dMuMdITszIOn1wPZPU03Iq/dQz9/6LB9/ClKo6iehgl9WXASyLIsGjE2WnvIM
xbccm34tPODNtYXYAFZyyiSrcFFr20eHxfoi2gZ3FhgMXtQVmXqiZBDAko+1/X+eLW6+W/U7cCXj
ZMSe3DK8aB5++SkR65EunX5eB0vcbwdzQZlKh2Vc2ycDVdnDGbQUvS8ubfJ73zPq4DrQxIZHuvUT
C8/7+vh5DLRSiY+rd+ZYIAvjykRN0s9SYsiqmXAqDu+EqkL85O7XO4eNbHXXU4a6XBi5B0bLIYdm
KDU2HE+uco873QAlFCVLLWsTFg+AiUIWt3BanncTpyZKtIGgHrSbmF4hBOb5LmpuNC8+xbFGIyxq
cNc8G1vgl3FasYg+IxlrRkDv9G5/AQupB7L0KYzJFybxxmEMsYm9qNd45j4htOJdIMuYjEcxnBqg
wHJTPe5jzk7kk3D5N04oAiqwZaiJxD1FvHNNg06w8vHeoeQVieDTKRGJYPekGujZq90Ufia68KJT
oA70XqPyiK14uFE7UIBd3ZL4Lv/t2cdgh8F4PR/Qgqx7t6qxCVQNkVmsD8crYXDJfcP/EXOuwerp
XHYFDyrOObSf82O4SMHJiDEUYd0o0AkZDowrvbHHKmMnGqW4N9+JZt79VoUSOw6/7l0vA5LLNOsg
20VbJ5fS3bGY11Ad0y+Syi1AeteAy//RJmb2AHBP8P4w3C9Gh+Txp0/q3JPmCHv2xj0x9BuO4IUp
KnRqoteJ379lcePuB8hx9zGHxnidvvwosXuhsOeRqEL0t2hhmAqvtRHsYzoor2W674bbdmYmd16Q
haDHZktgMt+7dccsXMU6c/RpwtaTOr4fkyquR/7kKWUpRcvsV3OcCZLXeCa9nZ5T+YDDK2bGJ/hK
2WZWC9+PtvfNRZeRuSkcSCRGPDE495ur31xVKLMipF3jZcKgJueETpzxi4grDjFeRDZUsTSRU55v
hUUfjQYpTFsCo67eaR7XtgoNPFAk6jb9tJpIEZW1YxunIE1x7lIGad00+TqrJk92vVnMvciQvwno
HGn9slPs2A/hPsGyDr5akFherftD/lS85HxBpkAgZ3YjEfvKDJ2lIkIgifh4ZB/erj2K87iAxAtZ
ZPPfv9mAD3c8rsp8mZbZQ8PvlVAZDm0rjlUw0pa5l9X91xXeeWCfJE/2qLwdSe4SxyeZZs/mYsbC
gpknFl+xwIlVP5QSH4E/RsIB07+C0q8DkGn3G6Irlr/9CNxMQQAA0GmEBem7aUhRwWF45hWYOXI9
6CbDt8I9OV0csMKZw1wsXzMvcsXd76VoQ5ZMo9mRBqtneyejZx7O2sc2bbPLd2qITavnvM9OTirh
2g3CniEzvcs8W6Y26phVK1hT8rgV0IwCeYPTnBJGP69asMUnOLfcV3Vkt3Auhn7xjvtdAnY9V/vj
MvQhl0/RAPP3jMBIxUbVBHVtriAxQ8ffq5AfCFQtVgcJ1Dl6ui/1gj5nQAq7RwEjqurLTL/duKZq
3Scxq4kzJgDvrj2Jxt+UOKR8c2maAACPdBpVIo6Xqpiq76Yz6s84Ich7lybAg/ZZifSgv849JVY3
LyeDMnj/0frQajVTZ32WXrITprUQ4YRDnfCkJ/PTJ5XljvCsVDHNJsyUOcK3Aho7/x0CiuLPxghB
XLWqCMr0XOVgwecu46mtYMJXaO1ApK1d9ftDg0ZzYv/4aC0K6sGMHXKTVWdTt7yEcKXy1jLLtAz5
IcQ7RGgAG8bFVyFIWU6udR+5T6HsrVUtpwO7OQJQ4cBHLtteYoxq6ZuJUYji2XsYyv2gb5rOmxuq
nqZFXBYvnHHlBD+KL5ocwwzL2lLOMMi2TMR3BkQsz3lGEQn3r2pJIVYOxXiGFTaJCgRXuscAVJGs
treK4LCVLN38OhThwH6XMKwkQnohOe6Mfgvpq77sumIG+7I90L6P441Nyk2PSPnhoS/D9GGGQoGd
8nppHhGTiBB4e8ADSqsCc3r9VYeRpB96Xe3qkiOHCIqPQxh+b33ovN9w1wf4dKkGkVJMLYcD3kx4
fCRlgCE3K0Ce4lyjXzcK8J0GTFoGf904MxKlk+WMKcCrKgg7MkexPgdZOLquJzo7iVeLGDGPHzn+
iFVQ/F2zWdkY/QgL4oW6adOxwxZoimFRypUDwKieZu+3Gygygvo8guM9samO54CFydv166flyzBr
X8um4y/VvxehmlQop9x3CvWCOWtXsf6b67VKZdpHEIomxqnEb2DJGnSjoA5qqrkqkiOn2nalVM3h
A3BGTClSWFFNZDF8/eB6+uOca+gpSe8UYwYB1LnfFBsALUvoK+S6P04au0+M0GCO3/CmKDtQFE6N
EIfp8cGaKu08xBC4U7i78KpPqsdIGqZWKuyIw54alPJg639Tb5k0nQCEGxev3CE/9iaYtRbzKJNb
uPYkrOrEIly8ggE3cZEwWuyviBdQY6Cbr1OfrJTaKFt2F00FdkxJ1rZ2hnpHo+bIluy20MBz2XgW
AIlJxSpVRzPQa0Ya6eMKDRmAk9G4vUMKG5TD2lyuSPom7y7tlg4bgxAVF5LWkYoc18JxEF9zvrno
WjKO/gLnDMUGQhwTpwyBWVT58ik0aFDovf3GFPvhltFHq/CFWtwGHi8YxDSRlrCuixrV3ymksfdQ
iBU9+LPpiRyt5vUTsxFWeBfJ4mxN86vvPRaK4kB2S28SoRtmPU/xR78XsY2OB/k/NolsnwG3dAyi
1HkAugxhfRJCtRGL6COUjqWkMRXEVmzYZxoeVYgg+VrONkvaUmq+6sFPegvM8kfr6d8hLnb4BCxi
IhHPC4hwT9+45zxmm1RylEMwTqfebO3pTzst1z8H4XcpgAbAxtNEWCm+vwe2yUYsTiVJ1U0nP/6y
eieBSvnkmQPOFLr6bTXGFvQn/WOR9UQ5qgJOmQfoZo+GoVjGWsGy6Z0rreWB7Nd7R53izcE7AH42
dUfqfMiphhgh7QTXtguqG8IQgDj0YEvR3UCEoFZiW933iNkbpcoBZwNvhMFJuiM/j/Tl1aWmFdR9
n6bHiQQjZary1NhM/ZeMtdFT6NUnD+HNpJe8GCo3b6NMAbjJCHQnEMODD2IKgG0zss4J5YQBs/7v
Xo18AmJ8t0gYrfBYtaU4lfvgBRB5hPx0GwHtyWLe373u7ZkjoReQlaMHm+rUwW6HVA/zUNU0xXYT
cuY8DZySZsbVyun2T+77DtLqhuuA0xhSnB6d3HEYJcQb5uoBv3qo6Ry3AN8wNUjrvXxCEP85aFJV
KbogaP3WVSRVEoqSWmUne9sbwZm0bAq1dXRGAEQ5FXHh1KHzSPa0COPFSe+brh8sdY9CzwjEv0/B
ijcm8cL7Kxd9Uq2fChnbezaePE6ZRVDwir/lUU8Nhyglh/913EUxBgJOAcoeDefmWob7uG+gNeGN
3WSZ06hvUnKyvppQQ1vmxM/Z5aGy+2BlLs/9nQroOwxBUGjRpUJHf7vuqemZUiqXIszI7WupmxAQ
2Msv3Wm9J0Aap7rGRIe3WQsiKjT5YQVEnVK0Mw8t0ZxeIZ8Dzsz9BT7fazNONfH1WG+6HVL6LZ0V
EyiOPO8FJTvhR7EWyXE2mqzX17isRnQfugIylZApYplqoOf5sNnjMM8c43FQwE6t+gl6U676+2Ov
hHo91bWd35Bmkght47Oao2f0jmRL4zgEmTKd0ffxKDC8VgeHXXrCnkPWYCiWEut0dm81haOnDBBT
KbAppt6C+gjKneWDKuZeZdsOCUb+YR6pc+N1l7xNOtG+b2apz4hu0bhyQbjNJzlYVLhY0JopBWTo
1fE/4ZTnNVeK7j4A3X/rpIpQ8XEoTl9aTmvPp20PEtSTvfS8mMru6V5epjodBVt6fI2PuWoGfM3I
zTQum7afePcOj9OzeOFpEI094LoDTIW/3xD61MXHJb2yUJBrYLVAyn7zbNWuf0eXvyKzNM8i0YEM
IM0yvm1U8a9hZB+7p/78TbHYRU8/A5tO6bx2zbh2iASnEtWj+Yu6iJWI8+2+Yo1YazfSkno44V3b
tdV5af4yx8FK2AaTDeqU/1y8R4Vd1cInF0zZKgx42mkeCXIVCkf0ccgob/WYPPkSfdNtUXvcgd4Z
wEJuLYupXc5lN6Aui3yilf2nfPDcIm9E6f+f0FB6gruBDym8MN63czAo5EqRlaOjx2FNxcJd9/HA
rVSjNmhWJMsD4DQ3t+etzn3lg1Mox7YgBwAaT0VHD81nbbOdhZL1UweOXaI0R2Xz0AaomspnNCr4
YaDR+ff6dO1JnmDT8HIaNqG58DUO6Bsdj47m9hEoemHKQ8T0lun5ltwwYAMkhedU++USJWfpItI9
CxFmEH/x6sJAkr9CWRG0QbjjGTGMXrmh0j9b2tYg4IkPVOYcDH1TN/mv85RS/ISMlLPM9KFojzoN
8aX+c1Kr97a14GdbCNpWSJ65MjTOnmXqBXzPmPbF5xiqC/MZCEy/ta+2i5ZLkb4aQIBb0XwdmT0i
mRLi4qoQCGJVO8kJb8fUKVNir5L1qJIeH0o9acqOmXhMQbH76bVWR1SbP8RGgApBR5RR7cbHeTHD
Af6tCk1MN8ZGdnX+U5UYxcmS5bSjkDl6fY9WB9JrL5wX4BQ4Oq8yug5Jmt7/du42mITUhcpKB6N9
G9q3fCCL6rx4ezC2sziY5IO/4RC+6juMufPsyIEqdRckqYG/nB3neJegX4IHDv0g7npwWm2HrDzJ
dqIXQT7+R9P7F5T3O0LbMBbMg7Zc/C5kNfuukWjvQO99R2OCPOoS11Xja2opjVjmxdNbFsGgp0pj
M+R6sBYa2dqzwf8fGjuLF2GRktWA477h5c8RBEf49a1XbxdJdZM/ypEvxB/wFXmj+F6xtcA9n+2n
/k8SxKvFa5WdOmV879TodWD9TlNAK7IiiDYg4P+RpUOArmlNBmsLqKrg2qbpsDcnw7RDYrpDJpyF
NQouWPiLUs3+M/yb1SkuKrAKKBZGiTJ6Rd4xOCJ2JMM+di9a70nWwyCULc0WoGP9nxN/CW+Ur9U2
2HCUlyq1k77zhh52az1rz19Y7mGcRAg+Da4msDb1kxSJGe0ukNTod0AQ2jc4iEZlmVkzSrUlYZ+l
TqOZBGxidIgcyYE5yE6GKEyrjpLPjFAh6zyabq63hhzpm9dtu0LbwAGNi2BwJnV594oiemzVyssn
BUcnectBLRVY7RoOChiEzsttiitFuxUanYY/pNa7mNv0qWrvrVws5M0AZY1Z9wFAaDAoIlzth2Nq
LR7B+IUNyFXroUpEQ/rCHKyodMyuyEDV+yoAeF/3ykWQiSo+yXEmThryHHmWITeWQnAIy+K4CTg3
Sqe4H1kpM/FQIv6Nlyn33atqBTR8zqrJzenM5JNsBrCCnn5xBdpHv4u6wICndVdMjMtpq9ejlt1r
94fDb3/AHWL88mw5r/EF1eVt8niWcUROL87WK4gTJ6BOp2VKVS3o+jAj+9XHxSF8pD4vJp5aD+wJ
d+ee4Pzha1kJyWdWwCG//2XefZzNHAlsLiHkuEQT6C8vM/C5yfPOOB3uOyvaMnfZRV++sQ7QVLaE
lWNhRbTPcokv2/wJtSWgbY9b8Q4waiMSKhbWH6G3RZEAb7bU4lQBV2WHdUQLrlKVwMM6VOlKgrjE
BhbONoktvVEepz7dqsZkjOaMrE5TaZcUZ8n2Lz/7GycvRPqPZBhHm1gE6BtdORMND9AvwbNQpkOG
JKAkV0gA3MI9Eeh/+Sag1A5wOLyDXZCz/FbFDFFaq9pFPD6dXQ7Kb13N5EPUvg7ESTetdb2WmP6v
zaKRS7qqpWEDb0jSqapqG4bkwbsU2y6TQoTPMksoow2g7jTzwiQHq3rYXjnKkhoPqF3g6xz5dzsb
EfUpGip7fGq1ZnM2wTQREXqIfY9wdsPw6yEPWtU5igwkwZURgDXL0i/+sc7MaYoZDCPg3cJKqPC3
PsUz1uv47i4v1APmzwO/BtzQ/SYHxS5M/YTxWRcAUgLvnYJrPp32o/0XFp9HX0od+Pf5ijRzyyNp
zCBTTNIOYIqVEeueN/fysFKggSJKHJIgvi0mjeNXsia+kak85gKcqTCVE6Sx4Z6HNtURFHYjJDMc
MghwMS0zN2lV3tv6rdqFTAhgTnuzw0Vdzp661Vwghisemh0VzHyKY2nL2i5KHBMY2+Yf9IZddHeu
ZP4VxSc19ufUCH5GGee4miQWVhPzmQizY9c/h7X1o5xGiyg403bkEPxXuP4Dsn8qPTGXdHkfDP0R
CvsvMJW0vh0wG9EJ/LebDfWd5I4N6gz/kLBd9lqXW/PmEo+LSiBNhZj8QDHkeUnZPPsi2hpnTYN4
oJgdPwOiFHaJzfiOTK/MvoKOnphwseZUt+ijV6nSrtiNMqzhng+fj4Af2OxibGFFfJaicgpUExNW
KhRRL+kz2ZSM8h/n/fgz/riON74L/AC4fvpNdHaEum9C/g9jHYUtQaAByiv5LZHsHRU+6xhJP9g7
0H0u3QBfZBACfju+0gjI06yK2cvYaZFLC/wPkW2I1Xmjxl37NMzoXVhRspcQcANS8DWgh9e7tzei
baIaM9SQTeq7clhFNX8x6NcRrEMtQDccYdkgzzIkC+spvX9tkvtgYsHerap2IHXB9fqkDTtCaQCu
yzVDXHueDYfVVllFCOnB4A24BJN7i9i6dWSE01a271o0TalkTqwc2xw7qgyC15cCsvjd/UKBo6XU
ittJcqRYfaZPcae6ic/svsYIHTWmmwxb4wX+txtw1o7VLB0doXBcPqutHQgKhmp20JEj5xXOicci
7bOvuY2KjYJ+T3WBmSQGHwzUufHNjJV96Gl5qn80dU95pqczOiF9G3tixFBcGMcFzZZQpdm3grW7
dh5MsK3FJRxU0deOwIGgYqSI+6Icr0Ap36y8rUzNxIySu0xZi2A959u8YOzbbeAyHXkLwRto0WjI
JnNFRpYt5OwtOLqkXiHn8KALrIsV4qR++6pmptwTJKKnoXalW90+6Id0YTqWDNMQLyKPiFfgLoWa
i8deBRivnBoFFpcjZlrn8GJlYdSTBEmRCqc3MkazyMofXka/at0ddMioJWluV6GajakMYQaOZYXb
yrTvTgGDbmSi/zd/Wj2jKwDXLpr2/T47duicfJrmn8g3loPwUtyzXucF32IBuCR7nrcWp/ErfeaN
WjMzwRFnRwXZJldFkWada5ED+XmcyrFVe/RI8xY6erFWYjq4OPlv/uezCuj5Tl9PEwodyRHS7iZo
TZKpaZ0JTwZ0tczY4hTtl84hzUfgURmQjhoIbp5kj62oS+zQcZLDHwPQY4sRF5kc42ZmnszVX12g
4VK/jOZiQbgHR1NockJqh8MkfXI+t6oLt785HKXqEvfkd8gbs/vDjNHBvjJWt98Pzu5BmWqKfdho
ExKtU7bH/Xz7U+tMCkCYpyCBimZEdbE7GQDR6L7loHxxKUTsV7T7pYcEKdvKAsXiyg/TTviHSjqv
ByzGfx0yEM9AZThCKcJOP3jIMK6Ga9Mv6q231JIMEAY4WTyoA3DA+WQTHaGK90Ni+IbucGCo3h0g
cPzkGU7QmyNFYZbLJtzWIFZGeXzYT7tJyx6zI7OPLerTPEhtAuxBNEWe4FQbJnvqvygZQ9Gj93DU
tM3CdiUSNGcLI/1S9sDI/4B1qaxKH7z0MlzzgYIvQh65464tTnnplZqadhUtT/RXQJshisYpJY3y
DIziLMAkkj/lyje9hprqDvv833DVbXTJMRHfMsGxv0yRr4qUQg7lxLAkxwMb3wrC1PO0UCzzF8da
0Ut/Au6J1gOP6g9eg2IquJnvuGQOPidHduhO2D0UA8Lma4WDJLltQx4ry845NN7wRpfwRyk3/Sru
1C6Hth7rnpSCiKUTUrW5xZQsnfHU2rF65Tmf6R+0hS61+4juYWnXCYs/B4UMBxaeOkpWRaYWk9fQ
XPbyH009I+e3ya0wbcSSabwyYSIV4IKWfzy0NPTVDL+haZrQUbsj0OFsW18eP1BNf/XIb8WytTTG
/wH8JwQH79Kjby9v1bV1CCPh7SDJoyQlWNyJHVu5XWqQzBRghBnX50cTAkn+fWZ2CtNq2mg8L834
zEOlN9VsqRGS7qYhJ8qS3musKVMzcI56O4Cm3iLGfrkxBmiMlCUyVw6uRP3N75vZcdhFnN5u7CJZ
/dC7czjFg79OQ+l8bULZXTxZ7byVnaPA3qifiaFEEqs9ku3iBmqp2nqV8KgRtzP1fARP6oxshsHc
sT9in9AxS8O05UbPgyN+WsibMKIErpR6VghU8hbxT81uvGKihsajbFyLijd5e4UkcfyUO/mMSawf
rOE8CeHsoSdvn5E/yx3AoCZfNv/mqmni6fMKOssaN4/PqkD6UjJEWJ9HLxdIBFOlI9YlwSVmaLak
31Ox0UPbtzL6nQG5tJrIvwTQ9Hr45m8plvOuM4K12tbOZ9AoGkvgIxvDbz2zEd1v3PXyRNl5goFg
noR32IJDRvu32LKDYDdfNmAdQ0jx6NwkGddXkK2eGEfu+HEUCT6Na73auTfaVQkKezpZ12xbLT/S
0hZVkhVRSWQRhXsM4aUROVbp+BYkp5XQ5SMoXI63/gWeqhqhu16xGMk8q2DjQm0H1gGBTNlCaHhL
RbhtS5bhHaOGBwaK8IlQnuygOElrcwIK7xxqM2qecBqP7eo8oOBmyMb8D2eGTnngK1opVec211cQ
vkMZiMLobqcvtf+AJG+it1NYhESFcpKArmpd62wEoIFhChrTdijMiTBAHqr5+Pe2oJiXqwwOMSaT
2HYGDVcdBC4SPZDYHrMRkXA9ME5fd3pfU36clTpeK7CjNc7pe0md4gDYAx+hJlOzp6FtmjnFDHta
o3TTwDfF/E+gNcXMLZSUxoPwdT+RDCGDtdFWE+x2d9J2wc72jmLm3phX2ghIAIdp6B+URpr1STQd
c40xqo96cCV+Q/h8uccSo4YfGjKFcWeroMnzkVnlMu1OY9m2jMTmPr7jebkGT//DboAdQcdG7dBD
wczKDDXmahH9LnkNIqZWsPDVn1d9BEJXa0TFTmWw0bjfUWCQktvwr3XdlEVICsqu2cNllAdOHd++
jQ6+iX4rU+kRcoLWI9KlJ3ZtieZeAky8MYOc15Ciqlg48x3+Omw5hcXHvwJ1Vj0yQRUjcXezWnOe
n6JUnRxCFzlnH+KKTrc55psDWOeQ7sECTJwCU15fuyxJeMGRt72Ri2+KxuubIzXpk6v7vTfsFYvt
xFeiBKDStlJ+0g+IrHYJ4rA1kUNLv9DO0z7cwkTbqEmuSOseqKYCk7/mBSHwXRSNxcDiIQTLZdCG
18PFyrqL+MxJgmfJ5LSAFAtXtT5TWKE/Iwp6pN9pBD45G3BpeOHiaOOl+Xy6KkuWUsj7qCuot+W4
IEdOHQViRYLc2zVBWJzzuO6TYqOpcTiM8T7T1JtGqh19QSws0vWCrPKWTfS98XMNRndCNvRNBxuH
zU3/GKQ9dygDekkHsTYTSupgaXNU2z8EY4DOUifgwWxB+5QEnI3y45WPLqEYlNWuZ5nZSB6J/WxT
1taWVaDSg083JACIyYZgBKIEAKkrI6lY9LLH9JUmZh906Y4ZhkjlMvYIXp3UY7g/eLyZoAxP1IfL
YbUEEv4XP240wi4oiP5SCE1KoMNGpgbAxbICseyTOd2d0rGaFFqt+iihLT48l9cVcGVwBKtRr/5j
2XKTbJHx4bmZF3F4Nshr6CLCLtoEV/sj1Me8KGv5PCxRXRvkij59Qack+a/lbXQVYNs0/ddAlBhY
yT2MVXhYqCyC8kpBRt+qhAyEqShl7LxEalTZ0SzY1Qy+FhqKok0LK5Q7tzC4MTpm4nyRJ46nrB2T
4RsuB7vY75H+X7QgFLYa5tGeztBK3UgwgDtQSfiRT/kNLAwLVmERX/ubCc72Pfw+gxtkwVSZpK7Y
HFL+PmhyF+wXOYWijKYaPBmiKepyYELcfcmoD3C3RPyPoaXNVVkf/etH9twSiqDlIuowp/be5sHe
9FSv+EKPs2mNUBydURGQj4N/vbybnhQYFi0bZTgjkUaMYo/5JQJoa11tCSYpialmLvgn6hqQUDmF
QcBqBSwenPTqDlENZ1nnRAUVnmUjd/qdS3sPYKVpkM+O2BufVCYHSp+ywtK6HT5JElMIQlC+V08b
+z8ymk8aw3OsvTleCFv1RthkHzmBG1/hZFGjY/vo0a1bCOrzjSiovlHh5e4c38eYm+10/mF+uErh
jTC2Pw5cnHn74NKDW0oMDiNgE1kN1NsvKPcce9z6A1aTDqEAUYi/MGqdG0Rhi5jZuc2XTq0lzIpb
vlKlLqJor7LUd+2A9meQGPLefKhXN6M0817YPMEqELRSH22i75nMgVwz3oGLqOLIzsOO2/lpdGky
x6eWfse2fmqd3WOD/nXAtUsVgYl7yu0ZC0H1HoWPuDQh74vACZE0fRPJY3jcNQ+dqeljIsM2FXsq
TDEbCEVqN59pgioFksELlhAirZ15xqYWIxoTMd57RgDbjL+ibcIv3ULZcMAU/HzO4323gT9GaoGK
w5L8HsI8UT5RUiE+bDlKUUnv2l8NreWcOrZ2YXvRnLToqUVytS17FfwshtyWbMExsDPLKtxXQnFA
vamYK+TfYWrc9cE5BcjD3q2iKpCWo/pZlvIlCHY1rC8ZM8hW0VFfExv8oU2JEzATH0r+8H9b1brD
pds/WiWWJvLDWxDzsQf3n07bieraw2dtlOE0ICpbjyyE1EFvgr8mmg6LPTmq0NELzS8zGoOEgRIo
OnxsMp/lR+GB5h0u/nZdNm4Lh634RQ2Vbau5GL/GS3eqCIiLISlMLHcwOh1uhkJsB92E7LZp5bdg
1rckEXO5COOSi4A2NFL2fUUW9v+j9XH5aEmDouH9AtOz6cc4bYTrGJvjpfoxWnlRd9fWZ9xWveNU
AHu2P92Gq/SBH/saH0Uc7eQgdOAVmx6MiIAXQzgGlZFpFYfIqdMut8ZRYyL5LpyH9xbUP93g5RoO
WdYOaa6WaBx0Op7f3I/Gio4wY72bwUhQcSJrrRDS2mV2OoPCA+/z7+5OOjcRtgDaG8nJA4OZRwwN
e4IG062h63yX2ZkJ9Vw/DVObZPMWPzbOI3ANta8M6rweUck/kKUdDcGxTPESMPlli0oNaJYcOfiu
l6N755WNO4yW9IoR+UDC1PCiKMSDOL1qrmy8yWYfBYuZQ/X51V8+t4rOAaThncfkHJP1kbmTOX57
Nr3R61Z95U+0BIDW6Vf8rW5uCoR8h4/SrBJBfsfnDZsIrpkzgfoTMlgnT1PRBmjSFr4NeLUUmYzZ
9ej804CG2mScmG5A+SjYXusMoFGikPk+8OnE1X5oqDTRKgK1q9cBI2N2RMXj7QDiCgEop86KeceY
yNIKeRXob2MAM7hML6WhMZR/EhDqIvlbJYgaz5qc0BurJCejZM5HwyjijxZR066U/uzRpCHwAY0r
lB1TVaRxbVt8KGOqjzCTqWZPf1xERPU4eDN4+3NdENHNJeSs9y3ZNXsevuEaKqbBMlhLgrBuxBHj
xbXd4GGb6ruijt0dBMW9b69SJpztHM+4feS5q9z/Ie9YXikz7TI45nEh3J2dFpAq7BUOyvsqYJP0
ABAsPPNHUsy8fpdLGnbZdqGwf8b2JQMWWIAtKWpqefz3wgM7EcxAvuKR78zg3ksxQ1lNGX67u/7e
EYnY2reMbheUsz+1M3B864ZQgX4TAlpsCvH+i+Cj9wJMqQRzZ/jiclWw+ACeMSPD++MDr8Jz85We
X3jMmGXwiF5bS7TnmklwiF+QtGSJzvbDqf5zPAl1G5FLw/U4WvkfgJ9YHK/ExlSo57UAjhtSBoPr
4poYlcOhUjEqRG9WUvSdYtNL6rm0VDtizS1mo3VyqdD990YxGazU6VPbNBW8lU7q1AFHpwHjSJdS
smHLsVGHVitNcHPGotDQ7Qbts12f1ruXI9hjZ6roAYW0bT95xv/g5iG064lYKYX8aIRtbrgcwD0z
DpsoeS9bbrSQivFOzoAxqb6lqO86yhIGUsNE2bccgLfStCLcqmTj5ybbLX32OlJJZFuOXizLhb8a
Sb41j6T5tbYymz1N3z5ITCHXM9qq+TiKUKAfJxfJvFM0w57+BmYXOhrDNM5EvrVyW6h4etLwHVQQ
J3435VSpKWs5pQMFnUn8fEvz0wxEf++GbeSMh5oPLhSS1ab0KrgP58+3OF3EcD+1sdk4qHSGKlNv
LNhewFhXnYZbP5y2e7cs8xitUyDmihHMrXa4fZKc20tK/BXvTK90Cie3IVt7l+JLeJuhnxNWYNJZ
VzTUDS8Pg146JBmulIaGyRSTwEOgMeFT1C7fbY+GZEexdc/uDEp+oakCRswuWgRHK/ldMX7sZNdL
YiJRyu+Yk9poNKy1iryRBg2lBfrkCEtsYg2FhebShOhuroJxb5vJl4ouvbnhWAsiysG8HlNhejUL
Boadk5tRRsC8Rm6LBFJMZTeQvA2b+0zNvixMgkbBTBXkaRsy+FefWlz4PC7WzWtHLqjt7GzWyREM
osPasxaDn3Eec5HUJ5Za73PbR6f/XiqUCUcSIwgRGpZbMM5B5xyRlMGYoXIaBX12LWVu83t79VTe
X846/c1Rwg6ME+EWTRA/J38aYmU+sZ9dQxUOOuMnN+go3AbOwhrafAbOnKmvoFZ14CM7Pe5XT8tk
DX2Wc6v3NUQoX7FfWhfKMdy62laGh9PoCdFVGqbH8TwvBqyOfd9CwgIO72Z9ebw5ApV7kzfPWaY+
2HQiQo7R+bncLkELcouutJm1RXUFEQpUb+/zJ1/og5W5aoEDZMm4RhjKqOXA58ixi1TRmeE8rojk
j1UF0bNfQ7TBbXApx2vZwPu9GSsYvQ792rbQPpHqBhtHY/zxGRWB7O9a4kbKDJVQXd8IaIPNXGlS
rnx1KMETc+lcibIxQeYUJ1xBmNB3jgNzBV+9GceqtXL2rjvvvNQs0j37tcanVGn4FjXk/51ukLH0
tej6pBGwq90s6/+Zqbu4r2Z2zMj2IbnjCZV2oGcxxzr+qazabrukelpQplCperrMwpigSv7975cT
4xgFjQDbYkmx0O5DWPvGVFKwxhCYb+L91B7caR2vg1d30HOv4t4HqcDeP4EbL5dU31hy2lhJJZHY
f2WgJd3jiltv1a8kGAVEN6WjO9RfkeOXqRvj7SxloGMQY+FKBIVv2VDj8IAnOiELoCWFA754asib
fWp1Lq3BuMj4ffx/T2moOfh2dmTIhZ2yfbZ8cWOUre78Xrsg3T/AH/Sc3+V5WAh8B35882NJhfZQ
HQtZ9dBTFXPA2qCKYnnxiVnnjXHsWXRzcSUtkXYXaKpXpgHhPyAJF6uLQIiIwELwHh3x56AQRBjb
bobWymZ0JCAuApbBpL8fATalPQndmJv6ygr0A69u4o4do5riFrg+3tEcWJ3CIakQciflwCUOt60M
Mgo5fwjssAG6GCYwMhAM9TyEuetJIIua3AFK5HxdCSJwGJJyOOh9cWDnkxbNHbjxqBw9snfni2ML
fe0SmIsNten6PXPD4rJuQLJ/8c4FrvuivaIHpPrAJpH/1W5bUORoLWOIR2tRJS3tEZZb3UaZaBs9
+9XMieTS7TXFEgRPDbkQ56vwPYVIvjjoytpoEUEZ62wqa1R7ypV8+8SsmLnsJM1tP9ImQFe6a8cb
VO0aVDLNRuyujvEBwXCwvHBwhoSnh2s5KW1wG0KizwLna4NNskx+uL9Zq6BQnZyMoOs1ALpAZsgR
Yx0XMCWONhS82qA+ilp5Q+A6h8Nbh7ievDka/pxbPED9LWAVrX9j7+/E6aXStfJyne4cF5qlEzwN
gPo9H89L3DZhfZV/V3/3iqzahkdGA/dXQMPGlZR2zZmC44kglP3J9zB176o93fJFhOHZISh4gkEt
Sw3ko9RwBoFGcGns+wo7YtA84WG6dzNoFuzMYUvUChr9OHleR7hDm44HCmy7TMFnyZgU0SVeUncU
enuQJVjH6lJLF0wcScjaTQskfd2b42HCHEx8vPNTpK0o9LWRuo/M89DYueqFC26dfhh9v+6IrktF
6sfjRui3J4YRMUnRLQkpFVQn//eQC2EG+wtixNOrSo5x+OznkAsAoGMcjbzD7DYbql7vc2dG8Y4r
o0puMDHj+JzDA6H0ZwmkLdCZRqLq8HmU94UxdY4Zoh75jTqkoE4T+lLglO9I8yLLMEHZm2K3nVJt
/KxRLE6sBmyCI1X7wqP4yPTSInWGWXh+fP6Ddazpfi4fbGmypdLH2eJjGLg/jOeU26mG4I0r/uEQ
lHkVJkBfI2WYBlCZC0e50fKeSA2zZrPbq77JuWzDDHzEZVI/wA7VExZeMikF9Lda/8L4na1/1jjB
ACOInA4SxFWk2dENlPg2NGkrbTBsL4huvnMpmX90g1sPI5DkNTAA+C/tNBdRf7eAxNh6jfFKXh+e
FPuwN9Pk6J3Q1C+tB/jNQeJjJio7N4L+pOWS510DVDLdOuX76quZbtWQyO1wpwS1xrumF5EtuzdZ
7uqD1uIoS07TeCSx2eHZNawEuApt+LEfBqru5wuyjUqLINtKnThpMMnH+0bSIpuIdNN/ebJlauHo
tgxlYlfI67W++lfFNrFqM4az6vYz8PMg2dBA62sdoghI2hhm1mkxZO33luBBIhpgGVaz7PYM2/Js
pTJxO9tCjcnvTfk0wMpbaSEpo6Zc5AiqbZtEAv2p3NLZT6TCw36uNsBhlqbttMKkaodAPYcXIEOi
s2/eYmki0WvoxjUSA0sQ3Axa5pep0qe9kdAU5G4Bbx3bCQ8sRwPFANvt1EvAIkfJxhC8CrV7R9uX
SsYgW1MYhYIWNPwgg3y2o52DCZ0Wlb+1+1ij9p7M6jQkqRpCZ3x67TbEZeXPsD2IVZRCi5dRf0QP
Lq9adc5YY4shmoxjdTuvleQRFGRuKQq+ZZj3HkK01iAjtMtw0vFXldYTJJPe0SLO7Afg5e4BGnlr
Esj2CHvyM6mbBP0GGRCEcs8iWMR4fZC5BIoTfovFB4EEt4gBUEjZynkAU8eDk6bEhfrtR7Q0JbEe
syijl6hi2upqZTzFF/DsOp/kpLVahxbaMUSIpMj4nmRua4g3XdF8GQ3AiQAxasm1wrASH4U2I+sJ
FEMF2BIHXmPGy6Wq5lBWio/Q7NCF3ldfWSIBouGHiDM9kA9kUxyr3WaBxfhtt+Zwq+t9YWpR0Lgo
7Q9OR0btg8YpLIYxMofH7sBbB2zjutgwejjAsHyHTm9Jv8rNGCXRo1ZawDDsHoIB4yvBrjL5fDI1
W7vk0PTxwUfRmqzEkBHrM7Ps53i+OtxtgR64fW2agwTQYn/oHx/bb/EizqwkkHJX4i1gbWab4Gc0
hGzzOJdrfQ5/55TF4nt7C9n834WsYcyectrEfXEoSXrn7Yiis/WoI3m1gQSSBMdanoFJHrrZ0Rgf
S0VkgEwhRDSTZSbXtBjiX4Fy+cfSHhgDkN2R/Ogoo47mZ3Z1yPl0Ktq2KulQMhDAMBzKebEf7vQm
gqpERG33DIP7vafWMJjuKBuOilVpOnpHcQNI1svTI+RsVbrPe4+zotiT+Aek6diLfBlA3DPL/gDC
WNNdSX9ajikODACCTQ4sb4KWoFx+98gjUH6J3+b2GLrtN4hO/MBERM1HIKlF2frhG5kVwfqD/Enf
/bwF5j3yZJjqoShKi8ydqZp+HRX2aI3qhyUXINo7Qglm6gpQHL9cBtg6NgnvF8St4Id1NO7yFEbW
zTgBohSB+pfyGnzM7F9fTeTh9pb6arXyEQ5n5bv14XQFSbDdxM3pFwLnSV9yQXx4ps1x1XnwS8iQ
xy/k56tYouus40dSmGzau5+WOH9aevgvcfuXQ1aoOPjhc3uhHUWxjNgmQA1D0BMNDSmFF2UhDQEW
m1LW7w91QnLCVjgbD/nvUgeQzNsB07iQHv20ZeV7k7cdhg2UhS+9LTNP8QxC3d+QmqUTOjPoDkQA
I2zA246PJsuJXEUgC2jDn+stbS6QysHm52pyJB+evNAinii6Gj8CDm4MLll34nHmEIjg4xvEctC/
r8Tfz6nVhxw5WWEiIdc0N7pWEwOu9twM3iTJ1lXIP2rEuJLlGCUsz8pmIc5vXTDLddyJicaC+G1u
/22iErsJX+h2P/K90itSTvrDu8r6PN7ixCwZ2o6jtRsLkbETCuykYA0lZNTQec+pb4XnL70Tbtyt
lwtAvEV/a5Lr0aap7x2TYZjuNtyaMxc1oGlAY350arhDD/oT6OAXJqA9k4Q40rI4DcOXJHDPlvFp
VF4zUJMwryZnyzgZaMszTXvrU9jM9Yw2pYwOdMCsq1uTc9Q4CGBLTZaw3V34W4wGEwyR+WHvpE52
BB0vyFyh/rvKTHo0pHBGoumNLJeSvjckOoSCFiMMza12FdpjFdi8yvKbgW4wmfouOZ9cA2cg9sFv
etAbrK03KTjGoKFGS29tiC0Zy+nt3Am0oY7EdGBb/oa/EtUgiOB3sC8Dff7iXL0Zmk/8Kd+xZCo4
XAt3vFVVjTyPxkd52J+9ao9faqWNR5FvAN8XtBnelJNHZJIgQrMlARTmHt6LP1qjLrzyInebubZM
Hf0Ux1YGN4OKMHibn4erPkk8OnGXAltYAvAxykoPJtbJSh1FurKgSCu5BY8s7P2rO1U/ZmT7ngU/
TCwzEBhY58kdOU8Oin5jsvT4mbHmzSiAUCxof7TZGSGvralU3lxsFDuNUwwuefp4h52vf4EPgYWJ
Nu4wHZnT1pRprSiIkno2iyNlnP2RPcCwT+oUQvcH6piviMiRCMAnKCaDeinL1wVzKYdgWvGf9Smp
GMhoX78ueHEm/0JLPrI9bdQrlhhleq89UfxlKePiaAub+87Xr3Q2bOlLWnBKPvOsfWwg7wK0jJ8A
D4vJcLI96KPMq7zoSq7M9cOECGvmUhOBvpLzXxR6DaA1IedGJXJmcOaGgBhOE4/g1qVpF9zRoXSC
0c1s4EYte+BLnzaOoQpGOpVH3WQ3E8x5h258MJDmxMLpcbK3xxCZaQ6eJBIzSMn3Sptd0DLOLw5w
8xz/aWDn1wP1WABaYdW2352L9YJNpcmgGFSB2h8SFSnsa2DOnh95u9EdmfxRZfGmN94rlQzYo6VM
K8QnC6ZYscgrY6LIYW2dSxcWZ9eSB005YKZ4jp4u38MFlN43++u1AbentgyigJazWHNJrXG1EoOy
cPIwe7yYg52LxGGO3x1lMYjUO5x+CDUXMzWTvpY1h7cTc/NqzpYpsD2Mk6FP3sZzVT9adSVHHg/t
7qbz+esISxMfKeU2owCL2iAMwH0odmiVCzpvRpUjpmt+yCXabxbPr1SexeNCoBN+tlXoH3o6Fbdc
dh4x19icyAcscJIDQfmpNgTYB/JomVw/dwVkQ7BqP31lE/yUShhdBiCkZtSsEk+aA+ZUHbb5iiVB
OEi0EPTEdbmbrdlhV1ePERAjor+Tg+2FEZj/USl7ewLt2sQR6MXxlqbwqW3t4q303BWijOrPPM/b
K4NA3adsFkAEdK4BLjRZkYkkzpGThUKoIuYI+dBOXMoyXLfyebt8YZr+Oyr+Tanpgy+3WLJD8wnJ
23Akz1h5Wa3B16SICwXLPZgtxzymIVNREwdMw++BJsw7NrK4deDeai+n2saAZZAdQ2A1K9iUWvN4
3c0yOxuaWmeCkY1/S+0uGJGPOKa2KumFmBuPd5PR5lP2TJJSBedcekxGupJR4w7nYxGq2PpGYIRJ
Vklogcy8ExTCXh46RJHtIRgEliKAQUvTxxwMW+dx1mp1STZf5q47hKBkdSC4G/wkFLj1lRA3H+j7
6ZCVZ+7rKtLJhjXrJjAJBENobHQoJQtUkmJjRRq3uWOoAomKIowJgIJCJ/bK60obUPFe57kJSdQi
sHKIR+mYLzsMwlrohH8XlMdnW0vCTql059QXIohR7OgcV8C01ZzDpiEgwgnLqneElCPrK4kchhWh
6N3Y+bZlLiv4cJ6ZXZPrSP/Ys83BNYRaODqMjHKOlbpYdLzjK285r4YmEqrr2oxC18aqyHvOPzGh
hM4grqlmLgRxXb5uhnueOV4Z7I8Z6dTWdlVLMXa8BJaEKijxxmkVRGt3d+p/rlfAGpEKWqcFlRbj
YyWb8otJIc+drN0hItek6sZAA9dkcDONpjhOKONfZCFcgtKelUFRnJ0SIgvXTN5+1Fw7mDw46GiN
i6QmTSZ7hkUfL2YL9KRE0whZq7XBOyfGY+d8WajH1wWN2Yv9L+PPHTuJylymyoL97Dr8WmW+HdeD
pT01HZB0bcV6sqSwsB3JXmWA6sPYzhgolCNp6GLaDzZDOP65Z8PelsInjj3JS67KmKLlewYujOhY
neDVQcRKJr0sVIPeBRUY9156KI1Hg+2y2/9fpgYdQ2H23bYyJHkwjZKU2u/R46WII+EvDyKkEe+W
/MDT+GcVNS2a9r+ranmCyN96I/xuso7A/llC0Q0qywcn23h+hv53aV0Q08/ZHHqg7o9EcyTIFKtd
lwalLGj5EXUNE33c0//6Lxg9G/xvAPJKAq5QnR64WBeNTcCKY+11ZOK5lx7VBaCMUQPDzySPxQIH
gs2OLuM9AtQoNTwll8706kOegRstWtLrpIJ01CLRJLqZW3AQ0UTR2umLUtB5pSkkutHO8THXEIxt
7MKHIujxiGcmYRO82hcLof5i/0pnPkGqfEY4t2AVGVDRSNwH6GJWB5uvp0dUn8f4PAbiG59Wkiry
s8diJRfj5CBF7rRQi4CWbI6xvIce1Zt4t0ZAOHepFi0HkISCGSnAc7V4J/pcAxV/rn49Y26yteGY
ct1bpOFw9HHR1VGUHLhWUFxqI7UxPmWzAwkx7Q+M1/DK/r9tH1yqscqU79FcTqrDe8AQeEFJcmzE
WqeeOvZlX1fuk4c44xuVzcMm7doVsfutJSPa/t1puPqnNW4Z7iR2pECG01kZzJP7XKeYcQLakoGD
54c2BvNfbY5yRt8IrYMvlJI6+zvx3ayZk6OdfUgYyKjKJfpTeLZtNLzWzZC5B4kAUPvxVX96nVvP
BNChRFeJnZ/BAaIxyJGQ1Qg7EQ7SCuVoT5sBvDRlpuGInN3GeQ4y6vENOYO57rBJTKMc9S3CuwLh
jsgtLDSQI8Xh7kdjX/NoEWpR5UadM0VpvquwPO7emGkw6TaPO4cTsuan2Ea7p+94lAm8zrKBZ/fE
SWcvQUuxF3ANJBiWuVg72YuZ/nnAkyULBLYHo3Rujbr1OxlMx+2ANv4G7p5MaROm6+98fXTh21Ty
+okZp62DV3XkSpIz4fLNcOQz/P1zlSgim6P8AJbf+ysY+eRDbku7dERBd0p0BU7RGmey7/oP7x3x
X1kaoBvQcRF77NnZ2mXRZUyZFAfgoIecSTai9Ik0Mpui6uxs0HMWQrGuQPz81Bz0v0BDrbT3ea7V
oaqQ5CQcAHPE06itBXhvwmomSGSc0rYQUJOFR981K7/lQpqMjC7QrBLPqzxyYOCY+HkbH1qP5INX
JUvZo6QtvrztBDK2d233C/EBFzSFirTWJV173xUMvme18MEQy3EgLVVARWjR0MBrXxu1V3pxwVs/
FqXsXh8Ho3ur6eFBTSEelhwAD2mJKbHq7QHKar/PqkCsNcQiYuR3M09RPR/Uc3tgwfTCc7jf2hPg
bpdamA22z+pH+xuQ762B6/WX0TheLfltqRCZ6+kYiOFYlMyifCi/31idzovYQxnpKD8KLPozzSj+
FACexJpSLRzAi/CHedwb1ARB7NPCq1kcRU6z6q+kVn0Orcqp1t8OqbUnrno2G+eVm8CD6Npyh6T5
He7TXgIDBrY3R/1HwvQ8D6uU/fpUsdGJ5meB6KKMHHbphHG/aLa1Bg7bDCvVs94fIVNLZ8oaMMgK
WWh4f2WTvHTtyBQHP9ktVuMnGSarsDqQz8irKDthMHdsIMJgeGgaFXFIdX0FbT5Tgeb/eo5PCHFs
E2NTdlqePzX1vUHeGxzhlzBE/z/60fuV6iNHg3EM4eHCgQh1hvLVDZMMU6QGnna6otgK9exu6AtV
0hTfO5hvaBpx6vl/oHo0/xuhiLMNVZlnSpAGFAMoUYB8K2fcz/3tY78aNB44bjtdKGz3C+mFhCwK
HqtHy1VqHZXKRf8nlonntiYZtkgCyo6igyyN7KwjllevKgpSRUmho4XUMYq7fkpBqQZikJMIVJQC
njMj3ntymIMQVDjGN9Gl+Dj3Htx6o6cKrG2Bx080+3FfWPE2poQcGcnL/w1UH7v5FL1r+Gv/p5nI
2b0P66e1Xq7YTQIHDWba0Vfx4nZfVVWRp10+pw8q2rIfw75eNlFKKvJ16YWRfv8N2Cb89eY6NXWq
sz34nmFgx2Zr8uc8g9Mb+35kZWwV9UtUrW4zTt0Jw2Ywz7Rx3qRDj0WD+MIGLH3U6fnPxGFX8E9t
Lj0Xq4Honcf0u07PyAc19PtHoSQc/2iH5urnZCEwhSnB2LYPgnTL6jEsKHN9y+DSIlp3ZA6oboOZ
vTYDQucR89bXs6FJzzimQXE1oQbF0AlPQbiOh5e1TNgzGqsFIaeBx1O4CSfF72SX5mIIsxXPDY+U
MfZE8SfztnA9sg4S8XFgkNkyCM/8bs+iYOdHLaTR52RAPlidk54ralNcdtmdnAv0Sf6Lo3CJZ0v7
0yvlyarksveFrZ3idGT/qLZTdOeeio1hBY5qD3ROsG9XwgNhqoq4Pl2/VP8A7ubluxuVizyw+9fv
4hqR2cQ8B2oBJZP8rkBj+7SFKe46TUiBCzrtxW4KI5o2V07CKjRUkwNyzmZmW2vw1JTMIHS1IVCZ
vIaaWqy+EtsAahD93yFdTH9eEQIFrMGzwBLC9NulfDpnqBAcz+DjSI/Rbj56tX7pgunWuWwSRjg3
Y5Y0b6xysZyq2eJ3Z98jeh477wx71YAbcKURUHs6tTeiOhFnofQUHdMVprBQb/UhPN4eHRPxBx0q
rAxxFf1eGsgRkPzt8+sU7fvVD5YUUyOd4qk3DrHQUGTF4nV6MKyAx6XxATggGdmQw2deEz7Gao/e
7i9numv2ZNxUQbDwMDuX/6fkTGRUX3alYvL36EYqV9UWnDvmzKGkIMYBomMUUwRx6o9SFyuPdn27
oggGp5xrPrj5sC5wV0bqOrlaSdGk1wr5uoLCnktehPgLFkYEmA+/FmxHpGO2QkwERLCSDKBT+waE
NXfeThd0z5qClH80JKEmdvbb7TQaSOj7LwdQVuTlxfF5nCSnQ8fhBxuo01OBMCW+7EoeZorJEC91
+QpE5WOPhcc7wgVmg7qwRH+dQnlE2Z9ZOyahwvboxQIizfeXBPr3Qmz+CwOrpMRGU3+hcG2OduAF
5LyxbXeqpMUfLjyG3RT3ECytrLyMn+EHVUeTqRRlOYxwHoepEKPSqg4Vaz1L73TxAqJM/SEPEIn8
gIZg0RGwDN2TRX3I5re7OVS4GacCtjmj4jN3Hn9dIpdkEvVIrY9TGg26yFFiV/yYLv+MUT2BAGrH
GxQq3SmxDwMWp+YwmduPI22LUaRpChMIYZWOu2lKLNkC689SBrqR2Hj58oHaoq45bMa5/Ygp54dn
xt6iJCdbasihgTrGRAZ+NFjwah9/EXuu/HrpqZBmUydEcR1Adkr+ZkyY+OvwSyk6/D/uGsg9txe6
lL1kXlNlXplymxye122d2wzx7Zm1DXvW/Z0m0kHt+FtuI/pRLBzDFEIaGUwG2+yP+aurAGEKvhsd
3wLyBUzB+1OdHWT57/y/zOS7/vYLYgkX7PzlP/4vhWANzmrRdgML8wpcgNGWkjBV0zA8A+vogoKJ
98bvsJx1PZ4oSReVO9Ma/uifa8JixUtt3pa3BvLLT8Kwlbr4T3xlJ8i+OjcIRyPj4kEPtPqJ94Ay
KEn44FCLaLd0eSFsrTRq7lbbI30iCRXYNUK2RmO/zfjeWHXILQnTLNhtcGMcXMU5AE4XQI/90BjY
ISv6Z6bC4C0+0pm/wXz9UVeoaUZJlO1gewcZwdL2tqaYBjt4cxE8JBcPkWLNN/kCkEKRdGtwFh6l
Tvub6N2FF/TE/qXPI/vBZZ3jnjNit/gXZ96frqCVAt0LqiV+/+4OCpYUM55IsRugZyXx01JjDGHz
FKckXVaFmtGUiA8FMMQwHP9zsjlvobvmRI5zOOatmquqYes2Uc7QLivTIkZNNYeXmhivSM4It46u
GFxEmE+GMOVUWyJQz1dHRb5ux6CIiqLWc7LEdbI9pcbW2d4mD4dF2sHa2Me/mwuBZey1TKj/lM3b
mlxK5svwXYjWgwHQ9lBuJguQy+/8WOX7sjojkTZ9jyy1FXuZDCM3UEU1Ue9z6oAsxdKU+7sUjkKQ
Cl/GsFR/PqlaDMIiifijtUAikpuOguVHqKGWsUkZqm+UgPlZIAZppeTJHPYK6kwlo6SeMemfD1/q
iCWujpIq20B5wmfBIKZ/WJX43QVxCSAJ9tueVHbi/duj27V4HCZhNlTfUXIO/5SVH8Yqwwx9vFKk
D9VbiFwu5nNknA+kX5Y3bS+GWqERR75jRw7Nt/5kPpQkUhEcaJ7TVRWkYH1ZeCfpk7S1A/cryCZY
FXpTLcKFs31/Y0b/ex8lzoRsMJOU+K3jktvVXNZp42yR0ZF+u1LqWPQY2r6WPYBIw9gTrEtJO9KP
fU8prZm1NLSsdWtMNUOlbLy9ZDTQdIhhjTaxJMqgCcgXRanlsEZ8zseezJKZs3vVqOkMxJZoC2p1
6o9QWe8sHqcNbZcdyTtIJhvb5SUwgTbds7tPiljz4osQijOHwXf9eCZAwa3U3knZ+1yVhC6TeCRc
L/a63P+QxGz7xoEG5mEbONTzNhhYNv0xTXV3gv0R+BtmMOrcgV6DZw952HSc2wmhqfNC/07S30u8
Xv86j3RA0ZkzZu/8/Nba6IWTNLZk+K6+mBxy36wBETwJ84mj8ZDOCTmf4Um3heIPKgHmsgemmXlt
sNQu2UEJrwHF+ZfYRhxcwYcATpzpvIHNaDmvRfREL4Fwl/0kUtlGzutsl9kjpmMR28qpJn/S2vz8
ziCqC65lych76Vpefh1vSgInfiJI+QA16zCFwOb2pH6dufpzDOCj60qDhmXDGm6kaBlJO9GZGs+H
OysatopZpsRixan59QlFBIEL47SVfEl28WjsG637YyYdIQD6IEUmVez2q5OysaFbXgUJtyV3Qcp/
cvz9P5qJd5VoMKuGPDQ/4csKU3nDmmsb92lLkI8l2U5kMGDUQQyZvTfV0kUJieHuUL0DdLZSQ9TT
kqpOuDQsTvXdAQ5x3BePgTNL3lIWPrPQqrN/EZTJ9VSmFIsmrWR0SyUS7lxwDvelkHqnYiBNbYcq
fCVUTG2aIMXy8pDcU+ii8azTSnVSkchDj2qrv80zr+WGsIbQDx0YpWU9k24JNS7YQU6wlSwcDoco
o/u6cIgzKysLKHXunTt3onjfJZ4xraX2/6kYvXpm36uvM5eR/Qem2QcgrmRmU9vleKvpzZF2rrOo
4nBxWX8Jg4rzwbIvlG6bM+C07jRejNYQixa2Ezbm/dOK9ZUx8CiHdplVko+DqBI1cE5M+qjVQ8Vc
bT8HLWkt1QEWfT+BFDtCN/18uzE0Oi5lXxy64i/7oA6oyMEH9ovEPA6gb+FjUe6IrNqxq9TyFghH
YUPUhZNohAPQkoINOUX1uZOXl1/w/h4Y1wGQcMyo+dIje5xso5Z4wppR4PtBIBBkGvgdoF21xIwY
TqOzNRLbo6b1EOetoSwgY+U6ZHoBERhbTqP7/vurUqpotk/gafaBxAFz0dzkE6wmnu3lS01uBY2O
eYGyt0sI+4siFP5/MXasNRmAasH1tDs1ZmI/1TqMqVpiL49pbnEeTGEPMasZMNjcmBCL7IaaQ0pv
Czr+H5tIFwiRbwdepQmDAO4K2QgT1Fz0wc84UZFvEoTY74pZaiqNpgCNa0oknqegRNQOqwgb0p0S
NjMYYJqqP+luacoNh117rysg4sQLqF7tSjC3wZGgn0URTZp27RCVdLAeHhObTX49FkC0DQWuVaMh
btrz+lTNlKv754CPPu+FOJABB6axd7wyiksy/Hi/TT7CaJyNRAwbv770fFZRnH3r8MdYdx9qsTJ6
OMzoCL/6BPVcjaU1L3QyDE4fEH/4I+JQctyz7ZsyXbUDPOH2BFmURMRpPYzNJ8iyn7SbZS2Xi0cT
x2Onjd5YAKrrlbKBo6baxZTkRxdCCmOaNBhFn3S++Cr4DU+M3aUFDQzyg0nm4m9y1CsMceIfTgYq
hnKjgQRHbBqVqv1IRIvCCqd9Yj2CclPC7Ny88Y0KmfVOTrZ/zVHKL+OhHo4WKqAvfqHzr3ySUqMo
2668pXnIT8wL4wGRrcGpPaESOzG51kfbADKghd6QXllLsepDuQmlNecY7fSoR7wsquYaA6pvF6RT
4jIoDS0SJP4CYh4889KmVCDA9G0hQw0FMIcaSDMQDsvYn34BQzFW0+MqzaLUuhp75IO52tUJ2/J1
feGNxbYcP3AEd98xuZw1A3q9igufYhlsgRrHg9Ftw1/FTJBWMlvH8dzG1SWLVwRuhpk1QLYptjMJ
NRRifPS5MGhPWVe5IpAXmBIaabmeqTDA0jV4wdFTRpJTYnv3ta1mvEWb1F4pD76aBB7pel7kmhbi
JoZxnxwMtJY4D+qUfX5p3wUCSHLSrOUFUMupWqC1lsO4dXFGp6701oPxIAxHNz+V/L0PwOHtyeHn
TkKCW8/Al9ntBBYm1XmslMZ9JGuoK6EKUrwJHMkct8kf8mtZcpJNCN3fP6yhVVqSVyArEnkEdgPg
cJLyjXLfmkXjFGXwGcrJe+ZPgEzdwbGXYHc8FeBZmId1qIac/fepKBk+TwGlP9kb7vKo1NeUCBUi
JAKQKNJQ0ayvw37v7y1CcQwvqvDR0za+KfjAN+tciIFwFY9Rv0n8AA009xc4jY/3qmeXsthM7fMM
gNmexcsmDtdot6rQ3ob52ni+pgyeMRap2dwqQJrFCAlt3X4iB4Ocdt2lqXCAa+bn9uFV8bFD4LNC
cGCc51ZHxTUocAseTUPIVFJU1n+MFsNKNJYIvEKar7Q36YWajJaUhJE/XMFiSUzIpV6ul8XhVOZ0
SaJ+cLwXfcY433zHKXaLI/AarIJ1FjGo8azauSvjl2aj9cxzg0ZPai5xgAbGkPLgv9xjKxviaqvH
+neZS/NKyGkWgBzZZCr1z+fwKdGerMDV6wgXAd/6Lywa7/4cVP8jaYL6EuhkcOTW98OKffXznhUT
sHNu+ToMtNybZqVJMng24DJUvr9auA+eR9aaEIie8GVbM/FaPVrWwoPBC7Q+QJqZXQnqbh2EcZTn
Jjr7ZfuitRsWhh2928WIIIv9ag4vpmE5SukJRJUc89ajBGCMwPSdmXStAS6OaMIZqQlxO7D7g4U1
l4XeK2qValkwZ54Mu1gP1iUy0kfGZf2xvkDYzTrsKhV5IESeyz5dGOvpX/DZWMUTZVdcUYllWR53
fugmFWKGKvNfWoicvS7/FGOJACMIzSSdy97Im2kb3gvdcy1hi93fgZEoW3JNZgVID0Wkc/zVRNQx
Zrb1OX5TfGCgSlHwd54pPNBFdSUXsOnleDGghUBfP6NYAXYJSjNMJp1R6OO5rnI8KB/O3JUfAZ5u
QAD3CpwyKg0q/rVt7JG/a+m6CyzsG8tI4gICQvHsQ2Dr2AS5/exrWMcicqT+QTJLy9ZUGPGDYLrT
KYfIbcdb8rxywqPqoVeJOoHUNTeF2C4SIhXfFaJrw8qEjPyKGji1xzwOKHxh+zLoSSYlx/EcRBjE
7aB6iFocGYyozejugOnfxSgv80jffeaur0H9UWTe+L5vtRlnUoFa8+9IV8WEMQ+iIYz2k+j/XJ7i
+OYMLoMh2FDP8txAUsAInjP4wnyuOPm8s5nKsiYfOrhlpTThFqwKVf0GbVBTmQOazGEU1n8VV2Uk
MK+oEfvklYRNtcIWTrvXhCaHG7mEqVqVCiQ1TEvYWhST1b7ca1tU9NklmkAdbB/Hr/DZmYMqMgcR
PV/+2fLM1DlThp1pRb/iJThOJtwxEi3RJ9GLmmfAtnKFtEyopv6LYecFmfviUMwMAJF3ic26l8lk
4s5Wg6XwMGNlisDLcx5tTmHwbwUhUQ4ATCYB2JmE2eNdsuTK3vd6eXg6MOjQDzF7G94SIHF85St2
FvBUxoXJVIr3b2Ez7f1/TcQLDbsdn0kW/ZuRPXUVmIIOX3ElLgi7d4Er8prxFZzme0PnxqQS3Ez2
Ks8GwLP4E9pfB1vMGnYdTTT0RUAH1SaemCNWweBcEm/K9e5QIEfEbp+xPwdvLTdyts70PQebbwWR
787b3+SHHdCVEE2hZTaIEfyCb2rXcH9NyYo1bfmlRlk2434AG5DSxgJtBXlO2RBMdCV5fMdd7U7b
Dph+P/V5tk9AN6W6+rVUdNHMec1q5iSvaYzap5zz9TkdJ0fYH+4QIgFXD7x8BScMRGrL0H+LwWqp
Ecy+mKeqXVnpP165qpa4Pzci5MtaMV3+wCg+3H9n+EmglhCYowhloPRNdaen3QubYVmRbGVHvH7s
f8VnxVQG0QrDIi5egCaghX/8Jjeo+v1IY3zpbn+QpNv90bYNTJ3WUg8UXvHBea/pJwSQsLVpH9b9
h0J5y/5batFlgEKLqTzR2K/gj0r3dazPjaIT2X6Yl/m0eH+AOHhAIJ0JXqiLKGrsF59sypTupZoM
lYfTsd+U4UWJXtXs7bjJFjuoqhGDiHS8rS0eky78/6j5gYGolUrvKHOBsmJ8sEWV6Ewptg49fVeA
3Qsqg/mpiR7ySf+qbt3YJIXte4u1jKAUlzFnYaNJsSpZLZ0r5I3E3x7f4afldvHE6ZYRHw8YtGXO
NNI6LQdxJ14R9q+6SYuj799jT7RFhqmE52bqMEFgr4TOCywYcwub8GsbPjmCT4CeyRk9nzMVY7oR
zfJfmPi6uJFooVYVZVlCS/oQZwJTjmQ0+sPWN6r4j+8MGZJmxO4fG0wfcFylV3i5heEtOkLISgeP
2UbJlXeaIwj/SgqxKw9GaMMhR/dI+LDQ/Zwxpt+i1JaVpjwKjk5h1O2uYBfyrfkN0c0kxRzFpDWS
V01rcVCxHqtxLGT+e3TsX7G5zCRG5WliiR7x2j3PJnjjpElnAcvyOb35JQkfb+9WCPPl4n4ENQJb
6gvZ+ruNmCk0RD1aKR0VoE8xErlh1A15Ku2p1mAw1jeQo1FU62I2IEpMYPNCJkDLPXxNAnps/f6J
o5GI1NqbIjlwgqEbPxdXKzacPO1cmIwxXDRIGSyamcYdlMt9lEjcUQhGCFfovL3686VO0j+onlPp
IHMr6h/bkWfbMvvz5gwyva7tI+nl3vt+6H99wtC0QUp4ZmLylJXmLlr/RpT0wlW6GHuQol22wjsg
OGzJGE1ZJSXmSYM2xYACq25AwfLEpz+MEPXCL9bvmkgBtFlGeevKYCMHiozHHM9T6dZyYRLGQnSw
/B/qx6/MF29UdwbrCjOyccN6ELCupln4TWJIGHC243Wu9Ymo7SFCat+EK7pvkjccftzwPZdHoMho
V84y4GKVXItW56k8fwE2wd2GrVzyBAmODsb6VXJvmiCiNxXCC6LAV5zl7fuTP+z83ZOZ9eiZq/s7
NcV6HHGpSF+Gv0UytajniLPSNO3Q5SKwZwzvtyKUkBFW/DRI4ZQFxSrnHkzzzvGoNlKcRXqKqFgp
0B3x799RHxvGkoa0I1KUwuYWGtNXUVSHt+cJ7wQbEygfD8j6tu+/mj6en3oUhgxNWGXD1rQuGs3I
EpgCPxkQrBCjfpYcEnV2vWqfcpiPdLSWxRpg6EOeksK0jPyaBKLXvDyDrHlMUzMES7+DWHeCIl65
8Df8hpxYRR0Gyi73dviByeds46uhM2BhQru3c28+NFpaJnURDPT8R81IZsA+Oh5VAw/1+CgT6MTF
/4rzbsl5sQ6fvTuE2jAUMus9Qw+R6fBJeX3YsqzBOH1K2yY9DPmT7SaHZM06Qi53H6/939chOtqA
KpUb/bxKiBlHU51zxvpI/pQ73DWo7Hvt/11X7mlyjDg1hU/gkoOy69Eu8tDIGdzdc5pA/0cXa2Lf
e8s+1pYn+ywBD5k2PtyR9lR9a4sI6f/O1SWgmyI1BI4ol+JQykLyaI+1BPpt2sBtFDQnglHg5ffr
AkkXcWAxfiJkQwrQhgnU4xd4wfda+mbiFBEczbSM5N2PUp5SeeGLQ/mqkBNgA3KmOvoShkXjNcza
SJGXgBpL47ACk5zxAi1oBQTBnh3r0zh4kGVXTsudxWTWW+kGMbUFjOuZK5wiX3FVUKys5PeBlk0m
oL+z1QJqzcrkNk8UvI8zMACIDnfOlGVAcPy56TyHmkz3UX8WqBDxVRNqCF5/z0l2OudCeKvbZjtH
yI2oWr1VsjjOCdwr5GtfW1+plXtVYEfT1Kf8vBo9P1umq8xnr9McVJ4rjmqy9xIZc0yn9gMeye/M
Y/m1oYH7IutEn0HB6siQCagzZylz6+RcReEwtDUKXDAcRUcQOChUkf1NlVQVrB1LyXHuuqMafsEX
R5tlz6f5QHZ3LtJQFieFRO4rHm2+T9muMmiLZwgwwhcZzGcfp7N7ZSq3AaTPS12XDfWp/YJIMv7z
gVaLeF4bJOTiEk3ke7KvANRkQyngwg0W/QMjlazX5nqkiuWgV9kf7pF0wSzVIZMWTRq06yPg0Orv
tyPkTuZtjVTJhA0iXR52PHDUC1xAdBTC+yJj7MNm5ww3ZIPUjvH61NJe671/35u5b27lsiJgeYNL
3GkqZqoZQAclxyevqpMvPa/mV7vtFxCBu58VHXeL+e4CSuGlozSxnaKJ35RX/S8z6PenrevGt8Pe
roD7KPwbT1q5iFhMH3WkGpbyy+UBe/SZzEGdvGDebICBb8q1F8oN2q0YPBIM+CosYwwRgXsRDW4X
JykwWaFXVYA2/6HLZ6oMcLSi/v3xpMfkVfC7m6Bt+TBh0EGG8srwV/atv/5tzf11DTlIkTrZUNLJ
P/iQz05f4XSJO8PyYGXC1HJ8ZykDtK0xEzZUnpgAkv26AcUlmv4T8PKRJ08N2aikA1Ph8DNyJuT5
bgYnzoWA29KBtuOEH+G3yOsn0VFNAgCAhvYsyVCmQDeJ0YWMAm/LUy3uXDKU1Tf1sODA7GOehxP9
zFrUBJmW8zRzbI+FN2gOqCEXzunzo2VcE2LZETvXaecM8Zj2DP3K3Jy+Ra8qxgtZplvJf3YxufT5
oI95K9od5L3t+e29cgcZioJaALMM96QjTkOqTfHTTnn8VS1jEjNSjblLcQnFuooV5ffkdxO/x/BU
ZDTUklTfZhcsx2x3rGu7IeTRTmYKnafkut18xorRuvKDA/dTj+x7w5rfDDaQ4GCWO1OvxLGIfuv0
Mod+A4iDeiCh3ItXb4qBSC+MLozhtVXbBkmCZkoqwYTcpUnFERvacCajrF4e4CZf6YSgKcwJow+B
BucH2UpGVKt2UWUTfpUnLiku3AmlHJIxznC/ny8WBMlnDcEPwF9BKpj24hTywjS0bZRAeTn2hoju
TL09BKVJJAagkmmsNcnzyDpq/WVLOwhECiupigphNjh2cEe2j8+MeTXiZe4wvIYbRDErmG0eqLlC
YyKISe+eRlMHH6SKht/NThu3nlCmO43my+3rFsKfdomyVcE9VxJL4OJZ/L2XbpO6Wsd5k+W3fG+u
p2HhceW/A25cgta2cura2dq20/A3eBVTk0aFsYnzaw4QHces+xx7o1LXfakt2dRd9qlsgC67Sb1X
rqyRX73XhoIxkulXlac5L+I+kC+F4DWU9mKT42qfGgvv/Lk+cPoVBqIpL2wP9L2aBXQtmAlOIRON
BKAff98ZLao5twYzYsbqcdkaEdl9Yx83TJs0u7Hr4Ag5DPQWRKSoUODGSxBBRrg5+WYyzJlPRVnc
hGCGV2mGivc8RB+qrsa1NTuJsqUT1/CUjiQk/Xewvdk2+2t4vCjRwCpNLG/0PodJ7y5NktP6QGSw
YV7Zw5UzoO9mTjMTcp131Srl8eMv9lxXJC+iSoFJXaNwMU88NrMnHklJd89olWd3kXpOJ0xkHSYB
OyKLJgrrdk+yxWOK34ox1eGrULZV6fmpGpnNc+Z7SnpodBhBBJvgbzfSi6l7zfx2u0AkcXdE62NF
jhjkYHsoBmxgH1cEjYUZw9wZbFG1Ujq3VWHgXyqXFBexfn930DwSKZGWm8GFNQ1MWivKtWka8XV8
ynwci6jLAg2yP2u+zdZfnrBT4P+HI0NRht1DY8R//BfYc/iqIhPYfWya8CQaDVUgoSb9WiihSK0H
xUAeL8YhVuHBXL4hqu9vgpGqpzn/gjt5tbSFe4pE62jcmYHWPghZdWjqvcySVTwZpzE4y3wMjm80
IhOhYW6DnHpDaXd4LzqBzHCm1tSh4zAI786ztar7AYtx4QskX72FHgj6zDzV+P5RlZdNiOSAFyQB
TGEQrmHgx2Lo5198tZxbQVvl0YkJpkA8kq89q4XtmwB/Qqi56OA7Z8wivJ8UbRz/yNskppEBWnYo
7aYomc+wQJp27RAfCPXt+G1acOCNrvfRdcWm2UZxvZ3RuoqJvn1pFTl0I+wHz9KIp5YdUyZQ9ERN
344hQhTLjXTRfGU6uaVUOYWk+zqqxPMZhZ9uON/d6xNLHJGDFPB7+vk0cYz+Rvrr1oEvxUIWHo9E
wtXV+YnxNnU7wj7f4u+SGu1BGP2T+wuDOsJeWIPegtoxGm0XA4TNDTU7N8JuC/vs/MTzoZmGEXM4
4DYxds8SNznivP5Of93Jqyrywovigf314RNqLv8FOVpk4bbs2iai0tYbPoPpGNU+anUPiyauXUHb
Mgg07a6Ofl+OsW4R1u3cJnMaMtExiqCKALi0yKDxj8y7yDWZssV9JttJrVs+T+QnCfY8UDkUORn4
wRhwIcP2VbzPW110V5yscBaqcqOAViWrFbjGWEV1KnauzoaxmKCCOdVqwy68G2lUYtFbnOEhir/F
BrywrBL+TDU6h3ifXNrdJKBed2hpMwAUtdl44CMN7jB7sE1kJ58N+CFf1RX/8Vhksx6Q/z/9hjfj
e7NV3BLJ2quDn6w5Xu6SoMlvwLGkHXY2w0n9CItoZWKd3yn3VUp0yQrIIqSfKSEm0LvY11+Q8nXR
6OHa+W0mE1mwXPuMXT23w4iQa3s1RwMaD4UPoXNhjvXF5zSHKBybZ+wixLmVktIgf0efwH8ZDAH3
ttIMg7xgVbCjbnifJ1QOuHVtn5menGH0AymuU1s56ttXfxSeIjlVlmK/7YoHJOEMOw5B+eRxiTyB
X2f7cOVdWOAudFlHjXvHbPa7Fg5Ya5xaOwU9Ak8z4xzS6SOWr9eDnlrToYU6LH6/Kyk6F9Afj1ip
HPLDMKHuWCa9jEqE/Y33ByYAjdKpPxnRMz+eTehg73H2wMfXWElrLLYWlLUhbw3N6pUFaXxvUOep
8ucfFzy4XniWHbmFORJmMlNv67He9iBL8F6HFdcUfpKzw5y0YPq48VTjhAMfLICmGJzP/IvpQaUg
Eee8t5y38cTzMqGUXn5GbI7F88D0ajNtO3EfF2Xnr3KpyUagox9nLG0Q6HvSclcmKiyBMP6ZwMsP
vNJlZ/AXhlKCNxEuHoy1x7SPZHnXry1IfzR8r8mHZIwgLU0zBBMgmvnaGIQcWVw0s15741eFJabX
9mJ0E+NHbkmWZ661Y5goJSJdYWZT/hDD1dfZnxtkLKRbHB4PCvmL9Hr228duo5nCrlnjXXN0bX4V
d02NAb/lNrVO8Hl3sId0pN0QwQfiyBMuuyV9eNny5D3UVjVnVgZdV0tLfYVyXgafE7FcLHUZRWXQ
Ik+w/8OTbDlarObsewBHW/Q6UsDG2x8dfyWbQHFLqv4wPVIc27spFWf29wxDjuT5l6D2OnCy6oDz
JsW5Uwb+1UqgKS11JrF8CQ8wbZNNJrPBC/zguEaiinV18uLL6P15N501v6/v8LxSQnqmn8RA3pqT
2F0IaStlEN9q+XNql7DAHM8vsDVpEFjolfdk8/aZA9sOVFvUQLWYUT+O7ctk4jGMtHZRiR2PzjFm
IhgGE99HG78impPrwh7pmLbqQKEBBBxrvq9g/xW0QQRK5BBVGlZcwyoWKmm7fhl8ogVQS7gPS84B
76zjij5ZEPO3aCo3c45nNT6HgRlRXvnJ5VvQoAfOr8GvLegDlMa8kaE0aejfXQoJkvpCSXQNc9iF
t3IN9AonNDtPbjqJ4dOt+8OzzCOpaUJD/cqpefj4mUKOy+n7ZsqT2cgPp/KK053Pj+Hn7vtBPDd8
+kqCsq4a7IfNLWUeuUbAK5Xg5lYlaXVeRZLDY/B7cu82XXL3VCrYOAZgVVaWOJxdfqISqS01vdb9
+LVPsZjPo4ZXEAnukQVUQu+ZYTIkljf9fvqmnIPZA/cxct7+haK8i/bfUmnCyaBxSqOcw57gdEGT
1Aam6oZLJEEG9siO2dTCkRFtEHYsXdBWTkLmlN1J/BFyt7we1g0WqI5WDlxeqwafU6fU8j5skqLF
KsWAiRGMoivyEyKNxGMrH/R0wTP/br+Wt6FUqn1NEGLoi/f5aUITqRSfjw6xpBB1Gsz/RGvf3vrF
uqleeN1N7ZqYVFGQKr4eKwYBoKSS5+es8WzsfkKvDspMIi4MLhc8XA+l0kRqMBv/TwSlEkRyGiYS
EVXDYlnDVhB4pvhs1Ctg63WmF6NM3/JEIUBiOck2vQcE9s19gCH04pWn1DWi7jxkw4wHChE/DtbJ
JhCLO6d86kUz7vHp+K4DPdZi1uSM+w30YpQmXZXCq30kPjJzcDNpvrwrgZBoIufD9ZgxjW3hlwvA
ZtiAMFkVY7bsRiMdJjolP3q2Q1eKQzMHWZmfCSBlX7syrkKRAbDr1VU53nyMDTyBLWefbqf4tH6A
CsAzmRCAFAzJWxDDpuBBhR3VfNcvPBklPi0ypipKMah4YYK99pMonZhtZWwdieifgpcBBVl+JbXo
1Dl+u9i5HzJO77g6E8ayKfW2sPW8j/sOje4TAkJs6lP0undG8TTkkoua/zJl6OaydR8hVXcKxbVk
/P8ShtSYOZi+5eTOvd+7h8x0aW1d3bwHEfyiQVsBuzbAt7OWVqbJ9lVmE3YzFjaOfAdvj9sHmPf7
zwQwEsPtYp40vnegswyqeh4n/0jpD+EmrDsQCT6xhRkkqSM/0uCJ5mpG/BeWKcW5TVTJV0vOyX4L
15IOWlI8O8Oj5LT/F/K2nrldA2acqSI1iqwkmvi7gHzUBjmZSTuV4ZI2K9RPpdanRKqKKv3cHxG1
pVfax5kPXra6BRMoSu/TRDQ0pyi/PTtCvcSf5/YXgYLqPohIx9dyHX/XjXcDyq1ZW+9u8m/ngBTy
oa+v+4rEwiuNkSG1hpSeHt3oJsidEeVQpqf0yML0L9oCo+Hufk47IVixTTm6+qJp41stLXmOzeV/
Eve/stg43SqwggenJ0pJy16zuiI5E08SYzUxJFKWF4PbNb16HD2/PYViqYyD9ST4ZkvoDA2Tfsiu
dEmbRocDFFWRbxIddhxivFmX7REe2fHqh5sC7x2TY44n4CwTmLmSWk9Fmxbv1q2P/zkxnCMGcakV
6mhQeXSEE7vUdGbBaNCC7MSlAUkS1tmginmuvx9sG9J8h2diYScTyST5q+THSu4rKzpT2f8mZTKy
wK8Em+zP4hH8inxfDo3IL5Ghn0RRMgA+uuuTq4ccn9v6Wl8JUsWYnS/+MQrjMrVNiEl/m5rg64ac
DWTv1V2NbvMPBqzCKGQC4DvA5t0PciiypM0IG079Kp+oVUERFP15ZLuKoS2ukxHypZdw2n9JVEgi
cM88ogL2PcwlarbJr7FpiEa6h05Nyttv3DuZELVrcPN9Cq/hbv/Rz7giXr3Gxvu023DxqOs9L2UR
6sU2TZrIznlcbuD2QFInz2BuF7bIKBs85ia5J95bse/BafwGaF4OROvAPVtoEJLR0yi/whWEW73F
zIFe6yxgjqmiCdR5ce1cGbSvYW9ZhWbDik9eAiXOrsYViG2EI9eStqbWwYtGOMT/kG6a04B6s3jK
ESnvzkFZXZ13slBanctKJ2Cu7lZjGMktOubaZcgUBNlK7c5qEahnTarf20/+VyRc/VNU9xdpK+Dk
l6lgHogR4HyM6wZ++YQti/M96OyrQcmkYljdJhZpbV5wOqEZ++04GgQdHUF6zRpA5fq/IkM8ZRvd
TuxpIkWiQM0KSRpUmBUG/dmS2cjguW5ySmz4kWqtLQBkdL1XFUQG+yVXbdvKxLDbHSINP/czyWr3
jSDokDdkhGDlbQ0Wim7qfJpgJFzKuNHdLJ7GlooqJi+YoO5O/qVOJJWPPCYZK4HcJVyDaQHPwm2W
MafYKu01ZuiA5Iy4GVWMkyZtcHukjafk5gaMM4nwximnQz5IEHTjSwLOziD+WZ7zAjW1T+5lzsN4
EbyeSnRivIUxHGXdnU1Fg47egO7EVRihuf+sjS+lSg1hWSNxHmR9sQN7Dy3gF42VAgoukWzC/G/R
fegil3r6Z8ELixkl0GsHEp3uEy5LjJC5J/9W01oIAbWa0XqM2WEU91shj/SbU7AlVYUyG6lC4W+8
TBYrEFfDuLU/jzUiltRfDfSqpCdFMFwVTKAeXg1lD5ybGErl6TjQQvV7JrPN6fCSIpvRkUL1TFUx
LzakKkEt6FK5FTg0yld/8xgs5ltMHyPgU8/kCLHNi1bHtsVDItmVtagV6gyCuA/ILC1xuWCzqlfe
LC1RTmbLdkegBqEao+x61DsEtsri5DyXGELRf1bvbT7vmqJxHDBnimAtN402UHZJ5HoPrV5cz/NF
LdTNLqh1zKSy38Fc+il7lIESPxBV/HSDJtuKHs5Fk6WDztcU/Ms7V9WSiMci63S1/mUc3X+DH8VH
Y17+P84Bl06CkYXR2wjy4Yo1RXE0W4+WpEufbxGMulJPOrRsToU6sEyvaD4IZXMpl3mFCvjGwQOt
RXvChkK1a2V6QcrYipSWyUw1XlIAwqWTDbMLaT76lLxyR51nXRS9GGEFgObj1i6RLOTt9vJW3DCP
6QJ3sDDH/fRvnJ/k+s9N2vVLVL6blNVgBk7vgGORNwu6Z/YS0pOxW8FycxlPDFE+aBPwnAmuK9eT
nVRfvb8/gYRD/W+F1bKgp8r8mYC5O/+1H6OL6Gm7UOjCthKbxtwbhkyetgfIROSbmF6e4zkH4A9r
EI6oQzPJm2yC/R0uJ650Qpg0CqWwAU7gGvZt+9fJ9KOkE9HzvpHwauHGnhRs4tHMfV5x7hAzAhkC
y9xtpI25wHKl/wAiLrWaKaOoy+cyIPWjK7HxIhxyFbA3Der0PtaJ75Hw8p7/yoN8FsDyDAd75SkP
j9Xe43DI/EOlnkRU+SZo6M1UyY2tSj2zLl3jtnrH2qpE1MoECLBoo6WVMbvf6v/kPoqJaei9ZWsy
WTp1IElVvQjA9nyHKaWXZPZ92k+6ZLthxvH42P4xIF5r1bykymM8TGmjJfEk6JxptStEQvAxffFb
VdH5mjY4fq5QJ6J177+KsDbQ0TES+DO6GYlqHldXT3IZKM8fVe5ZhuCpjVws08ri7LsRaKQXNL+G
XRIToIwE8tBvFQ7HvyYYfTmiuByKs3e2tZnik//b3hFml8E7IUv+ZbcyKGbNgjK/C9ehKEwkAQU1
8Vzoo6RN8FgiQo8uvzBv3Mprr7aEQ/xO8puZqld7jN133+KTEkETp5V4bXEQ/zSuYCuD65Bldawe
/yLhBQtjtQJRGnuNEytDqK9JyGIYcs4xExtx8ej0uLB2QDNFpwUhcbIQ7pem1MkD+esVnyTZURfN
55NtrdU2qu+GxCRIVJzPAaouSCSABIVU3yd/hUOjcWgOx/PQrVLne0ThKajpT6dESB+fvIwtVlt/
rtYDrckP4g4ZbzbuSeu0h/1HEjr5u35tYlcn0uVjboxk1FIgk2K3BbSSCZbUOjqhptwdnDKulBYw
ohCCQdTVhOjhp9v1wTF4G4TFuMqCagSBoHvsAM2OIQkbxNuIR4dN7AkEJ9SfoS3PGQUbFfCerf6c
SeESoSxVIYCjNB1VcVaOw1t8amnYN8WMJlmyTAttT7uaYIY1hjSxc7sYcZPm4zUBctObSqSe6vga
iaVfhUfdfP5RZeCe+QyxPD4VZYm7FYTKhq1+Jr3BhjUmQIING93d6+4uYRAid17GFWE+k38OuEbL
KOxnSU+6ryEwSWiYt1WzDhNG+LR4E3fXUW7xOE3M8ahM0OkhKYt4c/tV8eYYd47f7z0FUPBjyFjd
ZINs7kVJKqEaxjSZVc3EhZ9aqGmIVVgVIUZUwOyM6fYxuaIFFWX8QYKTMykM2Byjg6DemihX353y
1GzcODKpvW6qY2eHN5h7Bi4+JIDsTc2r3kBj1pR+2cSXQUYRT3z9qDTCZKfH/ZAOR/wj47AUW0jM
NJFnXzaRGqnoCjnZlkwWfPHzTjWut24evgQdwTsKWGZ123kPvODxsTIxtrXqULXPyLv2xZpimpVo
trQqex5/h5NZUsfnPNtMB5GXAWkNN4SFxOOiIevXaG0a/gPL4xWnY82fdyR8GpmvwJiNPQ1wTg7i
sxloaXiCsCBhJJdQmWRCHP5JTgUdi3hX69OGRGtXC42EIz0lIRHZlUQxKNR87+uUf88yWkYl+ix8
snp4mv0zUGlfBFUQ2B837FLswKSCuBwZOw2yYfajrNjknbqqXj68KNWAL/z7BQBnEIdh4vLB5BSQ
DvQynKrvU0tCEnJXe/hh5RVd3X9wglc1YBOIFijT4U/7dSM4jUt2f3T49k05nxETCka0QaPvpFvg
AEvx0Hp+C0JDb/kxgk3Q7pewxqzvqtvgRkgFT0AkHjOq8Wxev26xD8+97Kt5OvS9JCfwUoC8eMJ/
exSFs0SrHn63W9V8ht8m4Xaq6UsOX0tXQtGC3OskOsKqNmCmbPplAj0fFqPzzMSbtCaO+/ARQID3
T9bA4GpWjaW1xLC2vUDV1J3B6hMByqTQzvI+DWuqgMDXNZEL1PMfO1BVR1eyYL8KDexmr5jxCsOS
43VTD1AzXw6KvHkBs56VcLzs8q0qFxoAoVQtnIGz6HCu9Qi2/AbmZ6tVPD8DqOWEU42XOL94TfXQ
2UelURm8qwinkhOoaTwG2rf8+3a3bZk9UIylljQkeJJL8KAFd1IIzbAwU86jvIz+PTDFpvDQPReg
UpMDvORZ6q033wzVe5XvqHaV7csP1jChS0ZsBvLZILIaWKsfzSuP4KKFg/80/Sz8EWFwwnTX4rdI
QELtFnNeyA2FPYBIZ2uCYuH12u+WelILAYPOxkzkW6ZA6btFW+uajRTUwq2TavyP2X77aVgtOQnF
UexDQUikZh4xUo4locUPaYR87xbkMwE8eUWlXNDupE3Q6PTPjG+sfO/s13pwHk0rQ59m2w810eiP
FBZWdZ0Xy4PPVJBL9nckHe1/7JHUwtyeivyGyna/LeZpMQFIfs5kBDcA7V+tL60l/6iK7IskJ9UU
F8x6qi976IrCFi4geVO3hLp7k1GMUaPG7jmROrEAQ1110P/3GEa3vbyA/z3JaxES54jehdqO5Wvr
//Z0Jn+5Fyem8kpBxMax0SrJVKGENUU+UCbAsi5AdvM7BkOpw8vIbdmtzFcNZeaOjo+k4A8ZKQQR
NGH2ChEKe4Ctl+R7ARfwfjdeNdyAmCR1tBxYCrKW6uHJPJEb9M54UpXhR7yVZdfCEru8Mh8UnSZA
5ufyyiMKu1PalFTvUOPJ4U7CPvoDMKhZdhGMJiKfPymh3Tdl+JyDb57AgcVIHGrpX0hT/Il6th99
i2+d6zhbcjzd0oxJWSbN4xlblsffNnvjmi/eDtb7S6IDWnANkw+2TVDMbxmJDuAOmJnea/Ji4yqF
lM+q4URdNRDtvCHHWO8BzhdUwvy8OF/BwGaM09XO++j6JjUTf+zMGxLqZ09Fbc7KPyM8SNuAEYNN
iKI46waRQIzw0qb3R32OKMwL+XQ0gSjp/nPQdh5Uo1wXoJSGC9zU4vUfTvic8SMXmHNEHuA4QHlf
ZSnjKLFc1dd2UKK0op+DttGTzjf8DO3J05+30cb0vcuhK7zx9ulzfwot/mAhWZDAfYdfrwIK5Zae
15sSouSYaMAZTPWqr5CivKJAJCpFBEUe2PPDIknQ3VCC4HS9CMiDMqzQ+XXa8pQTCIhZPnj9DqcB
8qnS2/VY692kqA9JSjD3rLqZKXK+r3ePjZCOjgKwsGWpa3gXitaJYaOCsILapUEc/X991MLovoIO
9FWsTeQpHk3cJfjFwNjxBqvUQPmc00T70OlJW1XI6vyo2aGPHNX2LYaXxw4zDzn9HIguuKMPzIJU
NOlPTe2nc4h8pW5OIMkLExGHIm0W4+dFH4+gjeJhsoxZ+nK5WVEuGmaIWRHEPZ8UoQJmCPBR3FIL
gLXTVksZM1zeB6GaYdN8YvVfjFJP+mpFqA9ZQEEkBQ7zZRevbxDFHUXEiK/ydIscGStOpqupVu1h
By5qd2B9lUqQ53eQKyhbX/X0DSBKlE98o8zmqo1gIXppmgb3l9ekKT8Y82c/m1NYQnXOZbwE+yMz
GRXqeWPoXJ83C29hi7ujPjpRuA+WdmN2TOjjdu51J5CrZvVcA6obwCwzK190Zh0RX9agyR0q/VBg
O3BNOhv9JYAG0Qvv5z8oT2oYDUX0s2dWGNJ2+Z/Em7oOvdC1rmC0FpKJHxL78OXM+Q3KlYdtAtan
O1nFGu42/OgtR09QQ35NqsTD35V2pgen+OdGvi7HZMQTmAXsGNTdPgem5fGQ7tt0KiUjWyTwfL8y
6QuybC4hCKGf6k1U0mGbZOL9oXIaZ0liNhP8war3fQA3fB3wVoPrSUtcGrwlmAPIWmF1yvzmAKQ0
5QEfJri4l1Uam/xYBXIQ/aWjtIVVxgyxNdoq/HqhD1M62BA1AEqSmC8Mv8OPbf4SdnLxUqJ9hc7R
ydGEHgsou1XIyNegaJtTLLh+qTlZaxOMkHD8gkxiECYZ0D4MBZzysxalzz7hm5m563jJqt8pelF0
U364Y+y3jQM68JE33nfLWxMFPFHu/yU45n7cY3IOHkAzxdsKuq2oUS7Jca27DoldnOquCXvyKjSy
LvffeiwK3R9VSFOn+4Bi6E3ARK+/poZsphLtk4L7gGvWZSbw40hhl/8oSXveJRRgPTwXPwexfUJu
m4IafYlwm+jALpgk9bJkfhHqOQ4fK5RMEWQvG80fgJu7Q5Bi27+c5vRIwSKixBQXtI0gJ2uYB7df
+6fTkqShxX1uQqag7UtASuduQzSI39zmbuHAoeZYcGhKZGlhmrYMXU3z55DYwhR2yD1bfn0xvwH7
02tEmAWeoC5TZAT7jVp3UVQsJmRDFJk/XMBedY4Y0mvZtMa0qc/JsK2G2bbH4RCqB7e2iRUGTWP2
/9auPxv5O/23bCrM/HuF52Z3GcomeUydyu6mkBSR1tWLUbEB2vf1cdCAGWNCbVTLnacsL0NKoF3B
d8GCymiyBwWqTXMMMS8blAazw+xWom+buEy/KtK1X5dWb/Sf49GuXNVSMcTG9bl8d3V4+GWPQNaB
tj0KP2uwLIj0YcD3TZKlwtrISYpybcq6YgOuHp1vnRuX5U0FrjehCFH7WpYiP2O53bcXLWpOgGMC
rkNWQ46MREV621Rwu5V2WIgir/R5Y5s3JJ7Mf0Lk8DEdF/DOL0ly6Rj1Wv4LcqjY+gka6IGI6kBI
1V6k7vd3a3zWwyjCR5D2vNACX/o/FkRPz18dByx8R7dMDRimBEBggZbzAbkymm6Is3kKeJWS2PgP
mFAa7dn5MAqGa3VoZZqlYgcxYWgfcaB3XUoXPBsD9fqWfWunKnQ+VLsvKC85m25I0cPjzKAPiY0h
Mv547e7D/yK8CQnseO66M12uiArIQlsqN+cOQp9hs06a3R7Lt9huXnJJFIFlutGDrwigtFf7Sfcu
rYq4G8HY+SNENZb5G7sppfjdoou04+KcLx8otERPApkp+n/eAv3ocfS7ML+7crVN7hKWxHperaap
9rXhzuuD0hGzWEylRQXL7Jhd0piTe11BfrKZUEqNsX81ATxfGZmcbh+rai8T43DvXz0FlLe5AGSW
pVy+B482STCS9HlU3a9gtIgp95KqphTLdR2GXg0i9oNHbBh4xUFTodU0KUGEGwO8atKYROmNlgK6
8RFMFo81z3UdJNwbyA5zdxZa3Ow2s+JQH8R2z3jCNRzMU8y9/KIdXCU6N1X0523cLYpWQ1Skstxt
DQcRQoo43ER1w4onNjeXf5JKuPMDuEwbYBT908PEYX9AecNPRy4jRAH5g6zxok0LuYEWMlFk+ybD
oOaUkgEdj9bthKJtK4QFf6JfL2VJo5owDKGqXO52K6og2n8xNPeVCjtS9DC3ELBXkAvwNoVqJAkn
DM8YYq1PXB4atpDDhWtqc2HhkVBf1pdHrSzY7NRBt2xusGmyOCV3C2xfHmRY6uoxtUNa6ei+Ozbp
DjlaJmLU1z6CTvUvjwRfNj+04ipKUEhJxAiOYYA3GAvwsbg+SvUm8U2dIzOygI8vK3B0/IcwHzR7
DTbnpa9++CmQNksSSbGAk+Mt/ajDIRNcJIT45fKHLzKmTl8IxK++xqT8yeup7q5HFEc3KCDYpOiU
W/uAE3SEFOfS4xPtdWmkgcKLhPuV2DuD9RyqLtNRjIl/mkGxkp7TVApXiOmZEe3ICc7w4UHH1i4q
9BVeqwHhoCgphkiZgrCS006Hx1bf+qG6F2tp947taEkg81/CjNmaAilmSEczWVOWFzxb8SSDjyms
tfNYmx6y6tdZKEb9DnapG/d5Ysh0TWTQkTRHrpgc1k4Fzuz1G6kW/7YRRfDcX1519MokRYfeiHTA
jR2FaIWKFO7xygkMELoZwfkp5gI4W0vcR2XvyGpO03STE3ANhmZCCu9XsuVU2N/zIPnLbKezRqnW
Bi+YSuQ1F/QyS2mHg0PyfVvrkBydHTWORbxw9BRfc8QARls+Ncrf5TeSFGOQ1Os9VcQtbKBdn3RK
EFhMjSPhEsXWVMbAcdGw9CBZcFuZUPTc8VVenylZrXXLU4Dh8BlDitc7S7YvYdThv2SQw6tkz7CJ
QG60JUlH9WvUmi/w0h29ym0fV7hM4WrjFDqv+EFZzJ0ALQfFmNVz69sc6rbcPGJ+jGKKb3y2DFjw
//CDCrTIVQJTh8qYkF0e/UCdPyNVGxUAT6JwomR85uey6Hs++RW/XoZUnxamWGNitSr85/LCjWgi
4K9UBikaip3hp2BesWifJamo+6i4NoXbufp8gUtk2AXeUQh4PgelH6A/u+Jih7n6y+s7IqDGpO0V
drWLuqEzLwqrdCznFzHeLGyYP/nIN+CQp78sutCID7pp5m3UmbIJHSPH7xl5RV/t+pzVLBJDo4dx
PKwTVKvUMch4LUOri9u4UBS5BwUmutI0Km8sQu/kJo69Cirwz88sdm3zwdXOotsIwJ61h8K4xH1O
La7fwmZawilYMHMkwre/5ej/HimYL8necb0nyWo2bcJaer+kjjasYDoQdBRfKnF4F4Omu5VJMk3q
l671a3Eq26WE5HQUXsFGoFVmksGc5Vt19evlkYu9BHdcG/fFWKbWeVm5mT9tJmMSjtAJQWayifrg
NCot/Jv9zZ39Zotp/SUTyRno34T8jzI4ZmSVpEHb/h+kHWdNqqMcE3S7pd9bqWETiztLQJTRnddz
tnsyN+/q+0F+YWJAWz99ELzNuPfJIrwS6SxI80vgT3sabBruF7NsrCvsJBIB1ApD2UdWtmkAAf5a
8J60+CbH/wlWyr0VPi+qL0qxYCVOO2ZfVakwgzAbxicXubT9+dfxVREbjUE036R+KdvpL9LytsKG
AgXMyPIsGIFbQFbhXDNbF9ldcp2YU+0gwoojhPAj47H2t9i5SZf+paUNduLXtbZilgQ2kHx7c1bn
e7PJs7I3jRak30a9eGs5vcaM9ZaZyotZ/iO+aaGxQLDAhWpDa379s5SsyXfs0kcECEfH+NKAjIhL
i1iM6aV91iKruyYFPxqvNl4D5CMJfs8u5v5SmrRLwuSMPb83IAtJ1mujVSbpDjWClpr8uPIcwuW/
RYojcr0e+vPiIomxCZS0gUj56BT7274YvB8ZO0F9dOIjeKTp4no2t1evP5R1Y40jy7iZ77s1wBwE
QDGYur5vJF9VOYuvqgTw9R/8VFlPx0XbqvnY86FPdrEpzzX08zh0b1N/fjURywzXom+9fT8w66nv
B2/x1GlqYQd4mtHI7wVZGwiO2QyRKFquPv1tcd+GyNgp/8Njeemd9u1Awamgv/fBJA5u3A7cKFqc
+3ktpEFkFh2IvSaDO8omVqW7xJ9bcx9je/69gmr4403B+MglIvxbkBuus0skR/JmHAB7sA/RQUn4
urvB+Bs6OEIm8+a/mIoIAaRukNG++K3rH85NM6baerf5yujxBYnVIOUGYkZ2wbFKhec7vXV1B0KH
WRiLH4sN3LsY34xc/z25ExqjRvsZN4tfo+vhuqG10YA3TWF/1wzIam07kSl3asTqZtnaG6sw7PU7
kmz0RhR1setGK/mxKfmRaiKxLVRJkvdFXFLxH52YRX/vxSLjjR9CODwazhrqw8ub2pZQOXlqoXCb
HZZis4I1o+GuDhrCUuPA/eQF8J3GL3ItoViSf/F5bkZqvcSi2CSqfEaTc4zD5MQKD2B/PpnTNQNT
t1P4dB/gf8eJfVhc6IzF2+fZF4rjQHe8z6WHEHEWoNopnOdly+bvSjO8lgKXmWchrQTQ7MNEp6Ol
ytVCryMy0TPD8NfjJgqasIRrVV2GNrq0Bd0gZ+aKSMel7fhrFWn4eqstU0O7D7AUN3bmOsEqvow9
TKsGpIqKeAUqgxxpuT/lGApw/Zgwv/eDMlLZfj4uBcLAew2S0mXnP90yTYY8TTgES9kVI9ZuzSZg
Mj+1AOaiov/AZ9W3e5TRbygAj79icxTHqJX8FqJFRo7A/ERWSzkmvnY0z2xgPdXd2/EnAqNEoe/m
WDZLgVKry8vnWyYmAFs3rUH+0P6vOTEokQs5X68QwiwNt2FC/9xxzxtOA6QBbx+OKiFXrYpIg9+d
LH9cHXDBxqLET9O0+ZNxPdmVM6v6Prd1Khc9oKwjaJZRaZatVdoNgrPYNEijokOmEdpvyHRBgZQk
fnvWXnffGR1W5zPUbO5j5OtmVGYauy0Wm4khdKwvrBr90/RvPv5mJ+qjYwWceu7Wdrl3ID5aCe3L
vyNP9wpw+kuT4eD81TSqsjX/8U9CeGGkDbYMiVePbrYVI6RLeD8h4/cdZooPAYpooWWmo/MG9NOq
MWtb5l7jflgS7WDYB5ilmOQ3AcPXaT+pz83bOpOrvdiqi8VCp575knsSSFvUyaoUARreRyzdQhbm
nDEwLCreU82Pd4+zrxSZ/mSLdbAR4HU/W3vS7ommJ13420Qtsf0fjpEurvP0/9jI69yhi0fTZToM
W7T9y/DFFcMsNPmZlDnc0WkVepZedmWgDRB8j8Eums3UjX8g7HtgC4WlaVcm+oBnPMl8hXOqvgSN
DjoRoNgVOANPz1jjhOOjJy2wyv8eturlmlxYP1qlNyba9GrwifTkvKaVawPcVueKhDpUX7Ck3Fbi
L3If6aaON4nsY3ttqIP9ZFosvgQRYsnqKYvUnaT9xxEfqRtzLjboW+pi8tTah6mRfPi0XOQ/qhQu
8E93wEXmnxZD4HFM8uul6jKMdhkZXUHFQkz8Mz51nTcH+Fyl94jNJl28za0Rs4yklhTMeTNQR/uA
htTiVscqI5OUIM06htLtJ32rs29FIvcQ/b630jnZqPDNEmvRY5un15JQxHWgv84qEPulF3JXq60B
Zr9Nqj4k/F7hmFCocn2HQ8Y0uTpF1R8hkgt0T/YQ5SUZX5CPMXhw1rp82R+XrQk99ZdrQ5AsvYma
XWkxD5rR/Km7VNgAkUSYn41HIBT0ZzBsM6jR0JFSwkHyKpp6qp1T1NLWoMvYMBOAtzofz3EmZL29
lj20nqp1o7/5vei8qFyWtdSRd5NRv3sl+90BcCbSv5kvGwD8FFxVTfrgXivioTG+48z3cnS1L2nW
Zp5/3xgi9JYK3fJBu7KYxAQyZbfAxgNNmFvgxMFX4+8zjZRK58klCTnW16FNoiubiimdOPDSI6ID
MQljslxdlwgZQ6IFTvLCQCr3krq6RfCnTelkIJtjcCf9FNSJ6qtcmpTu3oBYiT+27Xh/gobqX//O
P4b4fJPxVsA0f/k9utgKUHjLAnXq3GnOS7k+TfcKVcuj8OvjbPcZnWSXU1UI/sOIat3S7e2MZMks
DqJCOgMWHDPHVXO4r6NkwLSap0FDMI78l8SoxC7wMTQttW+0Ubb3Xmzoi9kIbAS3aufhqc0bEhGE
N57d2N49paft+pzdfKSogKGcr3OKAF3kVFo+A2l9o43msO19E/M27f1/2XInxPkF4ZvN0TN/DHJx
ifyNN/r7xtrQ2yKl2A3pl28ekRyMbf5wDGfJoRt3GMhZtBS2JSgr5k8TBqtmaFxPCXQO+cYJ81s4
zSAol2MmtuvkOeoHvIhI4IscBlIn/pBmM2G0nXWgf1mDf6F92XxdsSb8Qkc8ichoubYNpCLbR50+
84MoxUc2Oy+NJL9NRvzSOCK3fqOidtXURlqEFn/Aay4D40o/DzQcUnlgQ4+SdPQQRJvBE3qEFykG
ioXmpPAu6bSQvs1zVTPh5Y+7Zjzb9DneTbyug38mhPWVpN+89nZbBOflR/gJcW75lEQJfjDEPzzq
RmYmaP5hqyVTwt84Jf7dnMmSEIL+5lJk7bDajhCGeNAvWcFho9QRfW6ZOK8ncpEbXRFAIqiGbG60
nIsLucOxsJ+oINncSgGPqAEAacMEgewMvYMkZDhzTjGQvDIOLrky5fXL1QDs8tzHinOIysdg/Cca
Xc0hDndpgeWjNOiNzySiFhgOj29rIvoG/IYz4wVxwKkXEjweDx6AePDSJ9BJkblJmnJvUslT3A0S
LDulJpKxHG8ngsNc9j1YgvIZMRnRnWJbj0zXTqhhsGPPf3Cl/71U3QhsM1RLJowaBR4OkDQZeup6
KOMz3yftEVUMoqsnVmGlsTkncAeCkTldIfiuUKtkugKh0kdMzEstDQcERXeqhztE8+Z/ppkdnbva
0s6A3fkR7w1BxxxyFgCqe9bUUDQvMJv6agie6n8+3SB6r015qS7DK/BM2qSpxUZtQC9nE0Vufrv0
d87swZzGi9239AyAoUgzRnU6GWQaRe94QyCqFuaXDhxociqjtV9jd6DqRqx+JDqbv77CrGQZYSOu
U6j/JxKOvCgYvNPMr47GcVd/lXFfUzfKIBiRQyjp6K8ooNkauws49/rxBMHAlXR6++5S632tmCiU
P0mhXC7/fWxb0Hp5qsVczQeHqEgObSCZQ2N0OeZjSMyzVuRwVc/7YjV9utIzaKw72P1N2nQR0vG/
BqEDOfuyy8yWUO3VIrT841cnrqZKUazjVce+Iw5YLM1P87FdgACd0Dz07KbFcRxWK6PfQe0Bkjb1
11NDfZ3++QhFhbRROpyeI5q2hN/XwrLzmmI8kDcmdvoTE3v62zmiiUKsLV5hiAfyPj3Dj0++wQ26
StRJW5ovxw3wPRztCiAI2tb5z3AuTz92uTMwQ4oAMmKV0qkH1E9U9adilOOQSJiJh9anK0wnZijs
9qldfEJxizIgAumwvGM3W209pX7T53SMNzFDnOjnXAKfircYnuxXJltUNwNY31FIV7COBxSvRwMR
O5dqAddgiW4MKzSqAKXjlEf9p9MzYf66vPW+eGaoXEbS7ZptR5zGL2FpfaOBQRBm9sXUMi1bWDzz
OtS/Am+eK0X0GPLPGmhpgRFaTXAxVLEBqsbYh0oPHRzZFyFbOMnByoK6L55/LohiwtOU5I+VikN9
++fWK5z1gq+g1MMKF2TUYCB9TuOEcOEAVX87lZYOGzqZVKXBJ81RuAhBEhgnqjUUZudWPJd7sgm5
AtRDbm+jXf6Ir9sTKFjwl9/t3DiNlEb0vepX4ShPUPJZXCxnxENhsZpGXsCC3wTtmh/RTy3ikwZa
Af6yxt3fvYBwxFYaJHMwGdLCKLQPKBN2/UTngpZVqiM8gs3+zmrpZANbZr7DKwsu2hgVSmbILaVF
4fKzDnmUIThj+nge7/lJ19UJfM+d8CROEb2UFow28PCwqiGR6zvfe2rMUeuAVTes3zyo3WE9Ktih
Pp5TrJfAmgAkrmXwOiVpkcfrSuYv6vE7koZnEfIGWGF5A8GvNUdvKnsMDJJj4g3iQ6hdIi71shpO
Pp3/Yg9hLjLJoQpA6w6yos5+cFO0CCGoOllYK46KgtfJYSmNeD9UKR0HPhoAYXEzm0+GrrjlKM/7
QAfTee4Y2aGvf8j5f9sNtw80ezmqWTPz4TTzoos4Xie1pqvk+D9pw9sdq+dan+szG71HolwfzOrT
tdoGC48mQCos5N0EdpluWkKPsOLtFuE4xUywfp7lpEBu3VIGQBh8CpPiqRVnxu43gdDWOz0UIBV4
GIjDHOawNMuB2ih7LRFkeYx2XP1H3523FD+imiNjhNUS7sUSgS3OVGchg7HnOGKokdRaWKASmVag
/8K1xqk0hV8WTJ5ePT3TKLTLVMQ/M6wTxbRgqoL2ZtoE9lzGHUHar41qM3oeNG1FMKlmcKPdjx8A
u7y5r6RJyo8/8xKbwEPoYht8Ehf6NMXF7Q2GAI3H5uVAI8wc++S5giItonbntcA882HKicTRubvK
yVqa7UtLB2RH3joS2KWKA2z7c5PcjbOut47VgDaRiP9Qv9zePoef8QeiSN1C9kL600ZdKyqeWVse
Dr5l52cOg2fS6YsG8NkKxo1H8pEvYfFo4p+wjmAfvhK0pdKKHE0JjW/xD+MIdiiqLVLjkCIDkcpp
podputhGpvPyF968NoNRtXcM66xyrmuR7fKXaCDv99Q8F3e34PDPPD+Ijl6ntWtKCWZvo6zclRE/
L837Q9mZOD8umTbL5gWPnzPLzKWHESndLcWCZ8NdGp6NpfTNL595XkFOSZt+y55MKiDCpH3bUEPl
j2FRLgeAxtmqVyW0gx5VVNPVmTwYBXNzeBSUz88D4uun790Kb27Nd8GvYNyp2HFq+ZNbkmcCvpnw
ihkugw0bK+qT2HNjaT1erb5pmQqTAeV6sAi6/+46pe5wMaoXxrlBDtlJS3x7JpemX2O4PnSeolr2
VInMyUkuJ10whKElVv78u8fNWBNVoWT3/whXq5inc7oGqSy+XN5IPZM22qlNcIc3LzhgU84cl1QT
dMqmuRBdNFfvaLVKzhD8FRPbPRO8NqMUDlWsS1aKGWOFeIYktu6L9U8CfvOAI7DmFfM2BufxglkH
sCXUHFk9BmUT9+UswEAo1vwjs1GFbTDi/yR82pPZOJ27o1BBLPxRDaBKt6gDpxICgNbLpAXLTE78
/vuvuGwTJUxlYNYvkC5JmXf2bWakNnn3rbiQ00rlv6PUjylOBQwHJKaIq5I6llhUYJ4lsv4ZLox2
ngLell+hRMaa/shKtTA59rrxnkx80jdD9okaVQFdOznz0mBKLoEO7Wjm6HaXV0W78GDQ3aETc7+e
7qz5U1zBdH2OpkqorYpfcQ72ibn95JfNEy0C4de7s4VWrOOZ5usJmqdU8+PIIU4Thl5+9T8oablV
slgbT6M3gTJ/zD+3Etn4PhdjRwIiSVPgumWJksGB9fWf75eO4Jj01IP9rC8MV0Qy/i1IS69tbY95
CGC5bwp7htJDhsWePIzPfz3OjE3q/16ndEfM7QabVcMIxnlh1ReZWSVEf15V6n2/mbQ7dDPvnqHA
8pf3rTocqc6DNHw8amZv8x6+z30gD0kCTbftwiXFXJO6quSIV0L1CRnlXdXzcHKqxzrCTtPV/w6F
tHU/si5koUrbFNANNYDKG2/iwveFmFgfnSoqGvv4ZrVPgYhaGWAY8mhPWvWhuuhr3A4Uj/vEdK8R
fvxh/hq82kuT293sBgw6uAbiikQ4jHoFglWqvUIHryUdPEq3n3Ft2n4NzxONu/B9+T0BOPIyJpY2
CdxARvrFMZKVTAOa7TKpy77WLNiBj6x3i5qWppaMuCOSVDQWihG65EWDGptabSXOndy0iW9h5+TB
SgHoZbYylMUUmUJ4uSUXeBh678qHXP7cioAZECrQ/GQu3AVBNDFcq1N7lTx4gRPdFeENnfXbfPF5
akSe3+krf/uUWpo/52aTQulhT1cGnRnzrb2PK8sVK+ljbsfRi5sAvtNPVkrgYbzS1UbYeP00A/nX
+VdDd4F1A3Ey+trnGoPSyHgeEYU5FFVGRYvNImT4lCR+8L7T7JVPlNfgzaz/QKe0K2J4AIpsLPWL
uzVfYPcsAU+HRatDghCWI4UcyAcoOZJApxuXiUTWEUsexqkXeBSxtcem5MpRUgqQS7Dbv7HYa4pr
UUlHZCu/6ODueSFkdwf307o8AkLo9UKNWPeZt+KEGLHYPMGXD6Cg+nkKNGHAuEeEx3SSzznm5HXA
cEhxgzPo4+D7PkUY/PD4bPiwwnwpSuuSCop6rKS2E7vxu+E/vJ8XZwhIEx2Pr3ihPaJRto6oouEV
kiHpd8UawP0PTVqoeYCgWnwrq7oCkrX2zs6m9nTKT9r1nibwSIBtWMsW7wtKomYYq6gV5Pz6TPHZ
HlCwPMK2328r7e4hXtCQCi3tsSkcbYJ7m8nbOlvx/wrrUA3njiwPssJ61k9gSc8lOUCGKHBAajkJ
/FCxeRQnFlXaUW+i/U8FVwizuRpto5DKka2YtKFAUoDsc9RJV1BuTtOthzO/bKufXKJzfG66Tq/s
1xAsSFZZ8hgZkMS/KZWUXSwvKsLUY43lCeYpg/kiNke/th1Cup3SM3lLZlLLjn+723jktMksFeu0
H1/GD34kI5D//gJU6D1WpXwhGQKJWKBH/IuF6c3yeddJDTirSiOnD0uAG5IbM1nzMRIUkdMU8bFF
CkFa9xNrE8ESG6OIfPhwKvVNQksoH4Bqbe9RB8HOzseZ1+leCG1EVfU8m/kiMeFERDJUFuxZJUae
A1KYKSuWqk383RxqBUdIrrm39eOuApaS5z0hEMeKrbxI9kEThbHpdiAFIcEz1/mLeSG8CMZOXI2n
B2lmph1OTyQz0owKqxKGYvfGtG+D7F8S38ERpEsKD8XdsZGMDC2xGtMGMaXE+qnOe0ikm2hulIT+
L9Q0zdyYuEX0d7HHMSNjbQl0t/S3htjLgCBKBUXJv/SwGE8MWOIvOUrE2PLYh3FhXsB959KvFwj3
EKc8vGC9CpS9XKVqnC9XaQcbhuHv8msrGXVDVW3u9XBaOgvBVNhuWCeddVq2BhVeoxuFsgTQp0nN
mnb7KtQajStEwKjPPrw0rMYpN47f2Fs7FIpsGEHEvdkHHsBiYYDH+o1ExdObq6Nx8/3XQ3oKL/O7
jYDSZ/6g1CDLH659x6qtsnlvsiskA0rnAkBoLa/QMGW1ZnrqgqOAr/VQa3fCVgDg46qGkDKC0C7U
VoUZaY+ysru8TtFZF9EoFqPOJxNIvb4VIJXftkx3OJgmE+unCTQhpzsx3J1xInPH93pld1Xnxc71
trPX4PcBQXXUaTNs054qoT4jVk7QGbbbv1BiH+80lr9QoqRFWM07aLTnZdJhxLxMxmIcmqa2be0z
xRCJsLeIIwzgQkqETlaFUOU3ELV3AznpOB7eHx7Ed0wPGZ5vGJTchkIdnrNvJpp2QpR967dEP4uV
Hqd0elkbdyZjiNhgNDy8Z+qz9XspX4ZxBk3fyaQI10NupVBUj3MO/A1MXSSEbTWGE7OF9DSKFwN5
5G7yCfn9pjGQ2sd1PA0GgXCSJFZCW+BI0Bj8cwCslDSXirfSFTkVf32Gt4xWjneFYeJMrSTeee1t
z9PMFe9wLLzAKA99tMHhXmfAiL3BuWZY/Dltgx+V/4a2bH+5ZOXNEMllcgUbAFllbkhN+P0juemv
PvFAvAv0ZqJr+Mbfc5aWKOD+AtJ+5dzmlWrzbiysGEQxjdF/3dLnWqm3ueVUMGKOZ6m3/FK+/rvc
mn86GGs0PcxTe30lxKAli0pan+s048eg8eY7Tc/tvoBqnmGjiqmnvpoH2+XExx0VSm38jy8OoANf
K4ZTYEK5ZZpQbQAiIyH4fAuldVLGrZZy4DQZQU0bYSHN8sKyNHFuZIBPGYx/DB1mDwD2RKwlw2xo
knEZrlD15zz8lQEqgRodcIWtp3fD+zOawyCyDbq9PmJ9f+RFMCzeag+MOpiCIcti++QhJTJWAOm5
Ik5wQPZ1QapZmS7Iqq99f5kQ70lQXEqQu2CQTRPz7xhrSwJAGa0sN08GMUnoc23igf5lyYaFCCNA
jFU8tk0hDQFruLmlENT3Xz/PlytrtoOpeeQJ1fgh+ZnxmdEk5pr9yPIZIMB5/5/JpT+PWPtynxYO
baSmrLZFt4utHIqcmws9gEtaxIEKrgJSnBHzWAQgXDN5xJzsD1vhtiLR9UQDPKj4nS4lPgfKOxkN
3sWLUiSo18yH3yhRwqBjj/Plvz+jOK8Tyth3z+HSDPgf0TKlzpqTNk/4Awm2I7CVXSrphnJGQIxf
/yvM+WGMfCVGOCTcMC5605VKZ2rTx/xhUl+NT8GW08r0OASsHS9QDgvHsv70n4Lfmmg+2VZCkq2z
7yvHbAxVMIJDfSXTQ2QAZovYExPLIZMYV2oldy3zCtBBgym11LJi+VNEZkj5BDc3eG1UI80RBxhU
6/F9Jra8q5IZvC4bKlGppBI3pjig8H2oBfgqB1YTvCavaIxPiURH0ap0EAvjgLKEWE89ua3jt6ay
Q96jTOXYAvzRTnhcJvXyuwqw/fRoDZwkCGmnxeQj7S9P6QwKu6cXazxrfNLvOVpZCS49U0vhXNgm
IxcE/JpkW+XmohAFfDFcKDS35UnXX6phfTsExTt6kEPHnOQPaLgFtehHwxv/QlLBAR2zsw0pDEar
mmjf2svwAX3+BlAcoQryk9DyeDiIfqOqYRHob60cgJpBIiyC37mjmbui7zVan+eZ6z19jDgdHdP+
ybDRmUzRB7bc47N41B6NuJwM45+npa/jHFTpCa6pRutk47VunoY/fw1Q8tBGu5V/G3uAXTqEaJbp
FkAwCgf/JnFYoaQR8W45+QnMzhKPgnM50WdR4r7WJwpxM3c9Rk138/MWC48f0KQ0ou9FhOeuRNJM
pAU7WSd2ecR5jC5efkBz40wWpIAugxJa8RMzKEQsHbj+qaYqjNlyzSxKnMfoTQWqKvTsoWhtWBSB
gQMbD/nZ8WZmYEPj7sIJUkw+6eaRqQIX6iQrsyAgscchl5up5a1NSUyrDr6JDCStoW9sCPQCT4Zm
pnq9ZEhcJmBAiSq+n+F8psIYHrQQ/M5tQ4rcELcLammG72/Uuo+xQa7FCDM5DI3xv0t/10FYqN3/
wm47CgMRfWnb6tikBJ5k/bPSD6j0US7Lkyet4hBCNaeyMBovU+WtHtgstxl+engz9IjiJuvzsAfw
oRIluYgirKuNt1K9RhF/hbJrHBJbgl9wdnwj7WuUQCKFCR8KLXrk8WTd9N+Y3cpVATzhHgICMUu4
BN08fqnUuOPMDt9cYlQXA4/a4RjJjMsqJGB6EAAh0+ALUzGeKaKQt1SNSKD6wwZEvf54HdGFuUwS
AMQHlB8O2taFhQzJBYhtXZMw/ZOUvFqI32i35QvJ4neFq0vg8gDEaL77KhUsac3GLkQSmnqiJynU
3Ma0l0vH2zMAcPy6uuJc7Z2ZSTyn/9jfptmkLPKnKw8y/LtmbS4PUfxUD7qkJKOmyXjz3sGfhroU
sa8Ky1eejkkVtyDYU7lHSWxp8S17ElcRqG3//H5QJISljSlWTPOPfWYMp7RHNtFvZ1zboiNbrHt5
EoqHLAkGl1Opr0HugIoI4wJTApkRRuN1XNO3kLtgTCrKWjHljWa0++iMWEFMbtPU5F9aNkbIIzjH
vzPiUnU4VPDSUGJ3M6AIiOPu/1imKStissQHKwO8T+Brvjkml3nnEicTjYPkJEd5bwK7uAuPRamO
X8+he1M/Ag2hbT1Go8+MinolhL86AYu73xq3DzNqdWku09bOwKqvass89Zu/RxSYVr9n2rk7IGIE
9t4j0djR5lpyujk+pK4wmcKyt1UAXj9lEJ6sKB0VnQ6YmPSL1PSVN8GhH9FqAl3O4oayOBMFKYRh
wpzxbGKzmov7B/A8FcHoA8sXjHbLyJ/vLgpKAbSVR0y9vnjyGZUpLVDdJw6xsS4vOGCh0N07p8E3
qp4SYLurEr0hXQ1ja4jM1l2ktW54dWlTZ6/D2SPU0dye/0ZiJtFjFLovEszQE0zJzcFshYZwp4lm
PFlSv5kY2q8Lh9QbLO8dVvuRhTb7gclKOy5HUNMQcOPYHBtOza6dd/Y1QRM1YaP1szl8t1UCrgoB
aCBpKQgMcTbmSiq8rPnaIVlyFrCNpTveLbf1Ph+9vbf8kEF4ii9200fsiC7vSlp6SqRc9TuDSBid
XG80Uml74B84k2cACp9LB7SbRfUWWzUI35RwARnbEvq5SqrfLsjAzeCzsObdasm0nJtjc4zL9Z/q
fR5bvEDT9pDiharGJ0htCEzUzDfonkRfNW6RBFXqTIQ4YWbg7bfc0DsKKI3R6r1PA2cnZrmRo52m
R63mRB9y18wMcQWUUG2LJrai11Zly8jHZO4/pldANXMTf4vn5tsy2DEpsE5Pl/e26OHxfqzZjU2c
26jZGLx0BXB0Q/Fc0G4L5ag0CqU562ZmZw5HaR8RtNzZM4dBEQE41hZIKK5jePsdG4i1fxOD/1zl
slWIyW6Al4AwB/gLg3q7SoMwgNpCgkJfhPK2AGeisTOoeQ7+aifN795UTinI2D8GKWsu/pXwA4+V
QaE/8/vkrOj97kZOr3+iuIwf5lQ2zBvhlFcI+U2rGbz+cE7+pdwfDFeGMSexX01XfrJtSGzY0+F+
x0YkxXsdtt0+Fvp0szL7zBjsi8xs/Bz9PoKyEfSgvYhlEIkl7n0+fSTepifBQY4FtZiSqalwuABu
DzDo1OuOTGFNN4d5KsdJHDKFyQrvDnnoQRSFVmpZUm5HUPz6qVvLHH90HT0zotKKTiC+HI+Fcx80
ZVBS4CckLhGD6uziXgX6dxOR1yaxjYnwo/X2jG/hvC61uSx8ExLqc18TfR4et1xRo0uyE1P9L/0q
qvUnFoyuLbUNVoeGJkaQBr8avVsUFMVqMZy2fww73YWaJ9bZSWMQZXa45iFx4h6loBjMOquZenTL
1rgoQrCzhnV43XYE6X5WBpZKtScSpP6ErHmeTdeffN/DBm5nTiM+yNB28tZGC45V36n9RtQBpX0Z
QMW1fCPT/b7EPetNmJa3jKsFiqa6GYXZ2qjBcLf0Zm/b5IKXoqoDmGzmlPqOhdTZEQ62pW4ZFxFB
w8bgrYUfLZd1CGnPDDo8GWWZ3iTZPNvphdIslKtqELPHfjH54Djkwsuv/Ekv8B/LuS+2Ymuk6usc
WbafCd8iYfcBMcWHaYjx+asgRF2HdxO7pzNOuPZLWqGd52sR/6vSJWCMsLsJcOhQrn5bdpkVyJ6y
Nd1UVbuk7COEb5b0cg9SwF3xJJRJL4B8a0CcnJaRf1kI2Gs8HL8kGQHJbQn+n3Ys0Y6ZOU+pABoG
ER1jvRMyR/jGTp0Y+qAfL2/XW9TID4TkbOrvxPtDTFcqadADkbP1uy62jKX14ElGismogr23nKC4
pd/73H9db7HMY2OIERJakvHOmmm1AgfLB3D6Bv4MrS4BzfEJQ9841nNHqmvVu5wjbV8hsFe/hh1V
sFTiyE/D7X2IxgVYO7fk7nCnR8AGrL0WHxFZ5TBWJnx0QYDBa/ydryD2obCT8oEVqFPSsYP4xGLK
tbm5WhAVsdb/ObLB5jgLxpWFutguO3+0DAvgetyHMGeANTtns64n3YNJ18uP+1JOMGJTsOs8g9ZO
Jm2ejUlgg8MvwnQXYHPmtTPnhj/3jb05J6ErFL0pMMLcFkOq1elppYuMXOQGbd5MMG4IjIB7sEBd
SLQxqjJxbBmc8YKtXRoXVL24vh43qkf8uT/Oj44eA1b+Wt0KvxiVBGRC+YPP3nOPOtbV5nMwFeoy
kUxj1uZx1YthWU9KmRd+QRxFn79TsBpF10m/fh/JOiZn9WN51ouvyN5VWhSMhEoSR4lg5IBPEeNF
wuDE8TmnuFLCsWqW2mFX50SJqIbolu1nSgGX+RwjprA1nWoSjJswfKqs4b0vxN5tAMF0YK0ze2ba
JhJ9NFek9mvdnVF+l0LjAmeaqVX2i395bCiLSlibC6D8rdV9TbPf7D9JkRozfE+h7fLKU5vrK8/2
CbS3eyy1uPH2zo6t6aEUhcnmdiBkqSA0fP1/Go6i9AzIrolED99UlSkNpLHk2pn29Tms/bHNzpOs
56bNfKc20IAUCizE25Cs69b2hQkX8pcTREiryddS7yAFI6eT5wpmHIfFZbLHW6l3Pfru6Tv8r46C
jcacRmDeptVU/jybp9plrM6osgVE2mh9M5MPR1maEPMkXQwKl6G2Pmd2FFt8bVpskidZbzKp9dOL
FptZO7/JZCgoqdL9jE2v0mCpqTTQQpuLVQ4g3+jGAS+887P82GDdqvroFhpSa0AWcHZZKOwRUq1C
1WSI+EXHIeZNnRxXDUJbKpUIwrmWCCKMoWB3lRK7oYfeZHRS999v7j/0oYEAoBNYPEd6pUDcXAZM
hlXTpmSZJj+AZWoBtOZ6FPIZqqTMVSCWNNJmApbppBKZ5zCR4165S73J6NYoKVwZnXvzEss7O7oJ
3FqQNcOrqXSS45y4vmYfGS16UHGHGWBvd2wED4QHmaV+7dnapt3BdW2q4tZ1br2IxFJpVl/N019z
AJMoiAr79Qc8HjX6JmMnCv3BUDW6wezOOdM1AdQ/8zHf8TpoUOLZL32uVoe2aLbe2d+4eTfcmvtn
6cqIDpk6kzEF0rBDewg0SB4OABj4QlTi6Hk0TlagwNOXth/eZRs9xb1Oj7Svu+ulO5p9U63qtYuc
lsj6+4E7JXi0CMaKiGZpvG1nYXWEYkenOk90sYUf0ZtBfFP6Q1W1/5gFJS3Rvc84JHO5E7o8RLgT
l73UckzyJuIp9mmNTYdKM2g0hezyxsrwPd4tuGkOgcA621AkPw1epUD6Hga/mKPqxoe4VUYb2oAX
AoSkVS+Gl/blW6jCe3+c4BCWNd/ttkhvCKmx3x6Ignr6GxSPabxVINjvS7t+UdZ3fQHdziAuSQor
XHEkwM7VCn4G0KzHHsU6c0T1yxAQa5uUG3luRkKwhpbFoCh/IOjif/cLAlXUvl+CUphYLoi7P0Pd
qp5EMlX/OQxs7KECx8MiX7oXhEJXibq3n5dTIDwzvM9eja7EYyg8v8a/6A9EznMinJKIBiKLwY3g
ZCwkTbRlfwmCZDC1z7G7Fj9rVWKOp9ZjE+FkH3Heu9qVy2V0sZ6asg/9QE9zyPRewaHNq7zHchQh
mH8gI7qPUj2c//aNVU2rEj06Q2yvVtqhCB9jbp7nD5/Rpwi8bAmIznDSu6Fn9em/4bSQNDHhIj+m
gO4plBU56zi07p1G8AolKPEh+wpYt2Vvro/4INsP9FczDd0NPX0jUEkSbK6jOEHlGTBvQeIe54Rx
EmBgJoV7pk/TywXNLz+ZnWZcgMGcXUIz4IGd+EvOvwSCe1XQPqb0RBZInzZIeZ5UgBqq6u2N68Y/
xU93RCjUtoikCbIReTbT8vgd8uXm1Fe3PXa6RG4NHS518b0WtyrIHch20KJT9s7N1hvNDn73k1xL
iPw9K/gNOqx4rt395PtOI2bHfnOE/SULbmtn7jGtd6jJ8fDiOvRXJn2ejEXk7zNdARl4yYw9eUZL
ILtNqlmWY2TjrtNen6ixB0i4oJGTRfPJL3SQiCbO0LQfavjqnOfcUUrdEtwjWIxB2MM8vSWwLoNS
9cjWvyR6DZJhe+61oMe/g5fr/ywYFMSKOICHQEh0H6ubp7GIVZVBDrdeLEAdFWrYD9fjTYcAKpCk
XGrKKJSMyJHpuxlrrMnrOne4O6c5jRG898rgatNlriKxJkUzR5nxtmNTmKYO1V6ARcoOx6l/4lA/
irB5VQLR/ZnJdZC4rdrRttMn1mu27IsmcVWebU6Vx1Kn7a4lblQllAWuOEWZwE2MmitiCdF6Eopv
df0qNMxy7FGgKfIyp9GNhtmfAobgRfl8W6CMEk4KJMn4NJ+XBVW0w9wBU2oEosxkKzs5wZ0SM26/
aSFyyLnN3jGiL/4Q1Vs5LPRRr8q24JMqrARqy597RYL4EWkcYy/BAObK5tuNrNNuAV+0t1Gn0vae
hqU1VMIR5oWmXV4FBAWNaUvKQH2vZWowbLVMP9SCv7gFt/4jkmwXfJtIVEBLr9EqT4xA7MEBH1Xe
ZyVt30EPJCiRa+PZk363woDliMdOwlGz0Cc7/WjzxvJuLrXp/XvktHvAGUMZp93NhI2eSGOVM5pG
iJPkieO84Ndc3wLS47ttWg8QmDhVY9f6jknAi2spbucG9Qr33evZuR4cu0TrPfjVoezIVmdaRtJ6
aPjExIk13M8kpJoGPF0cLDdPOI+kGzl6y7cgkzGTe7WvrDDnX2RMqlUxSm4JUg4zu/+lJfh+yi67
0BYBWK+UIzRHv8jrqO1XL8baWzBkPBCsHfhAepOqqfLMz8mL3HPw5750Wpqj/1oh10LcPnbZyBx9
sPvP7wPHJTOZnCOj87XT5MH/2LkJNYfgV1/L291S0ct5cZgbo8l1VnTfAFlNQ2tboY1tOpY1wKxL
hg3k0rvK7mRF7/x2EH7wY5QZgWJ1NzpTG2SNiNb7+VAjaUDmNDO6BwGq/Qjgy2EB0ggbrHldEGks
lkJk0LYIa8GtjANnIEKyhNU4y68ziie56rX8WyjtHX+y2jtHK0XQhmY7aCvjUn9mXzeUpfPOZNYd
Bq7YLYncyS1wacKleD1W63wdnVBpncwiHjnnttAanfzD0HzdGo6ZSPYj8h0+43IIFCAEuwQEVVzc
9aS+Zkpyz6kclmrBquuCznFoIlXzU5huuQgs4DcJtqdtg7b5pasnU30hsaW+1CfhZKsTFQJ43nHp
IC2ImE5szH3DG6vrCLHbzTPrX5hyY1tjtGsgpRtjx5eZKwDM+/G+rM8YL7a7Hk47mHE/Bp53KqJS
Uz1glq5FP2UhOpkcC8xwAPQIzdAjwgAVK9E1xPZKLwGf9e49ASQxKWbDNTUzBVDo154TKQXifng2
f/HkGfN/1EgIipM2aNE06atUE9N+X0+0k6IKvr9mlBCgQkt91vGBAjHHhWrsKcCTztQjTOVXioK/
f7OEEQrviB0VLRGGsKvOvFzdKbtDiruF7wMeCVNZLvMYLY2ywhltYGmYplxoE9moOMyxIMAXw0z7
njbngjDwu2SbM1Mfb8fLeZXjcZRZLt8iDAy4IPL1bTRM0T6cbKPphU8RQdRazdKOl675237lM5Uj
oRI3Jmu49b7zHhWFnyIC3dAgCBpd6eEO79PreAWu824A6a6N0XWOeWALceGotT9JILZjo1f2nb/T
syN88KvOq0bzd8Buoe9Zvs2MyVNoRjGmndTYBeXpZIz+dyk9rDjE2cqNjsYtrj+OKTSe7F1cVpv/
o6swduw85aNyxVQYzzxflSG7GtLzHM5uj6zyKmFhoHcJtrGVaZEuIT116pPp5oRO9LfQrCKdJquJ
AKilJIT2mWCVWpv7z3iub64fwUH9e1HKGPQqqGZL0ovGas1KglgqbjlrveeVyiWtukXpCfpUf1Iw
dv80IejdGrR3h6z3ZMZaOVhnI5SRSYpNbsraRfPgHMJlyQsMe03Tq6IO/OyHItTsqarGdkcyH0aj
ZnJqfvKMDYfEaANDQ0SshWxyzFYnjNEQWYe9Kf1tCbTeHitiUdvotcrWXcR+G18e83pu5dgTT6OT
pU1TID12pktZmAfDECiZ4FzRgC+v/+EJk8/aw8Vd2omF40QLPtbM3RcEJcvvQqkn7F06CvHH+g7i
Aud02GQ+8ffRw50KFilyGqg3gzTKNtHTVbBYTgjrI7CTEuDVEKoaFM8l4U/dd6S6bR9rVZxkoARx
eAAP/9z68+uRQeuCaSWHffxrrSGfLhvGnQTBV7UfiOML30tl2i0dZbFr3BpTzp+lkXK0T49FF8kj
tcCuj08063WhF/7qczLA0KKnL/ygffzVjawg/8zkBHko8QC+RnjTTCWqmVqv9ONzhxqnX68R1rgR
Dda9KJzFcaxJcV6fyJ4J8QB9zqebrCSKzX6nsMjE6MuktaSArRE6Mg4g1blZi5x26Y5+DEtcyOwf
pq6J9Vuvd3ZZDId+i62NYEkzb+Wh+kupdpkKUHcL5KJhS2flGPSH/OjovkPxq7aT4v96DYBa9UtR
ZiRdwLgDkWfT0yNrPUkg7XOvdlhQ5veBtET1lCmj8TLLG5wlMxROtWHVYu7TgSJ+GEqzdh2Aw//t
8jSLcEPbvD2E+Ub61jTZNay/MeDrolWuoC7iLcmZViv4wB5gXnUN7VJeP3DQ4Fv9tOkyg9TRtSh6
i5O1SUePF7cenz2Ag2v07teECoZrZTGmGqB+HeIcETjmRY5ip2suvBILdhVcdHOwJVfLE/zgmY5r
TsThz2w+rpEsTOYwXY3MQ+ZDzds9neLnOLnsac+q9/dBZitfkMWe6vwADog+BnNxc75YSJvD0B88
Z0EHUSuFdUVN7ddfpQ4+pmzAt/ehR4W0YCa34yr7mBkQxWqc6gn1+TuNZnL/f7BbCDpHIRlmp5+Z
YCD/tA+k3/EgubH0ZcDCiEPQ2tTGIPr1i1HF3DGfI9fO4lFzq9A5tqqbpXJT1eoIkmcYwa1rq9m4
BniWWSowJK/OOdJSvJGTOKKxGperezYFZVopv0j4voCN3uKdk6RjVY+FzelJi6Jzkli6jiZRfawg
g2lFG8UQy0kluRtKgOEomEQooPmSszSrZHEa7ucAui8u5/CIRLOkEcfLgxgEGFzIDj0EUtRcE7m6
w1XJ9LzW3Ee25p5CWIHdm7Dly4B6A2oN4iTpPAnfZFqKJD+hQIaO/FUtKSbqcMru6vAHQSdhftpO
efoVbMOGUv/tlgtgnsUmkWo3QzAWplSZdkPWaGjkwWx/EgBUj57jumQ+kq06X4dbvcAHMwFmB2Tz
S6AqNlHBC/K4YUyT2FUWfO6TwBB8ZP2PXxlBBblAJC89HaVnDdmQMupMYq2s2pUP3tqw9VnM3fK6
T+BedLyysCuanbeKOn11oOtxYKJgYF/+runzW1AKAxbyRO27nk/LIxrIGxtzsjl6cDiQBCuXyUhD
r3SfEpGO4rWmnUbrsgVY+i6YOCgXXKgBtDFbiFYWozuBDUXhi/6L3O1cPZ6TnfwNsICBjWg2aHPg
PDSqadu7ecsB1cWcUx0jQRot+20ZumWLpPX1EO90o0jkNmJ3ShyxQweTIPtJgqlr7StLDrHz5jlh
oZ8VHkz2kwpn9gpjJ815YAAFNXr/5HbAd4WVl33CezTImLCjchaf48WdfP/IYxLCAWKXEKpSta1n
HactPEceHMMsW+96tCq0u42ECJoYYRnmShIjSL79JJr3u8Bc5FV1xPXnf7JnZ1D71a9wd0E0Y39x
E1EaU62UEwbitSToN3wAezUxptNKZHijQbV2PUVCWgem90oGPErvJZ/B2gDnOCVs8yr2qDcTj+ZG
AlSVceM8iZBdcHei1qDH4vdguKC6pC6hxDk5i6Em2NF65mtMzPgXMfGvu6CqYwwac6DmjJkuKSSB
NxUSMFKcSYQpFZgpqd/he5eoWXFJh6XhzlNvhGjRiJEEeLaz0FOD7i2CmDRHw7uCvPEgGBTUVZJm
lvwFlqjIjSqiAOthVE7yqm2E8PPXOGHwvmUdW0lWozUIGdQ7MRlRRixbp9e5GInz0K8uH+l34+9H
7eyhsguzX0z/fHoJpISM3MjsNNyxQuYiwQwt55SiLfvrt4Xr6vnTAYvnz+kOZXjZc5Af9bQkCqTP
bCRWZ1L6W2A0TuGeva65h60UOEKh2RX2cLQQe/sn+wltakmx88TZFYF5sQJIv5vKzUp1DEam2u6k
qqZcgRslEIZMR0As4dYgqv40chzUWg3quIUTOfUT2/690Q54ypVaXHWoJS8iKCAwFsfBP/fSiTdA
8/wpqHjbYguCHBIOXcsz8yeDgjwIwmDYQt7r4tgFYg9QNhfa2LtehDkqJBP3WwHlHizmg86YF+jy
yxFEdX2H+OPfaSMdZ5adNWsDx+nzO5GNR2i7vJefbyjUIq13+xq4KIbIGC9JczOlViMu2dNYRzML
VAZvibXOlxobAQRY9v3121HG6CNNXdRZsMg6YF8P2hDHwsm8QjoLflW6WneDXQaj7VTx1Au8inf1
BtcGpLluFK7Valhtuid/ktkhYLi6B+WlQAghD0o8jFpP8f2lIURUTceo9LGKmLjhmUCBc8gYN0rf
sGSW+VS1b8ebcI7Qw5u9f0wqjPakSReoB806bGq4xwW/LymOoeY9HZ3z7pIcXUAwW7UZ4P0dy4cG
VM8iRnz8JiAFy196YhpKS0CDPuwob/X9nJxRHnq+HookzVOGydDnwJRBMPjMs/JpSaU6MUCvNqIS
WL6fCIiklqyqDErhMviVTYrOGSOGWokMMDGvuz5tW/6TB8Za249aTRW9IW2BvtkDp6k41fPMDkUc
nUuTXCmWsRecgd7IEPsm5HZh5cj75fuYKMwpU/oG3R3Eep4xqH9YH4KUYfnj5BELZbMnHGQkixWt
nzKJsw5BXxR3TL+q0X2PWZ1jiXwEdBAXZc9p7lFk+Hr11NiCftDGcCRlDhSUGG84+tju1DdJHP74
YexLijYn15nlK5pe4whPd9yLujMdQMPotnF9j+d6G4VgoD7wkLYTVvB7EUDVeCduIYfwBGQiilqB
9dgW9dIDAg3RagZTpJKf9s3sRA6j+6eSv5VH2CagNTyttJhmBvG9Uo7dCxCgdBLuIW3px6B9qF78
kA/HEWx8A7RV6XGnrdl52lYqe4I6L5+9bEeSm6EEEVJNN4tVGlK+Vzmbg61+w1F5KzvTfQ+sgs0s
wNZL9s9JBK5Nz88RgG6QC2yQ83gMeaonqR5ER4ar1+EfBLcpI1/UJVPlxIRT6COPpNEE683eXJ+8
1HlWNjIGuQCdQr+EZRVk91EnIRji3FsrD+M3ogKWRNfoS50a4EH8cZ2/NoByC7g21OIkjqx3T3Kp
1oYlFzc6T1BB9KEFIdh8FdQR+orLrXDUT2QX1wE8F7EghzzIPFJkVxCoODPVX/INOUtFL6JXjoyH
KQCbXia7Rmu1rs20PZgUAeIkYU3irUIA4ZCRiAUwFWRS3Wb8gPcaUXw9DNdSsoP4fiKT8VUa5hAO
4n1wbCPv5/RsTeFWH/SbTzYWWOfICQceD8GUyHOzQOuE2hOFtwyAqlaVKgdXm1TXZBMPmKuxj5SG
XGO+K1rdJeM3kJln1hyHNaK3VdVQMG+3Cxn1gXiHLvRk8gPKBz5+Ky5FCHyBC0OQJocZnQJknPSa
6pDd7u/Rb9phSzQ9RFLJpgMveje8QTxkGKMrudyz1kuGvVPj90dbLJg+7N2FmPLd6DDq5LgBHIhe
zH8G2+8vgrCMi3rG7bqazz9af4U/xKnT23kQJODmxnS1MBOWbSjShT0TEOE3qx06/Xz85RC1hb5U
iFEJSDozjUsEKjfmgmCk6O04LTVvh7lPXaZYhirfXWLrQD4vyHDLfd0+BLNPfJ+TBkFRPYBkQTbP
JFeC1OzNyAeUtJD53y8UklFEep8sEqKBsCYmBLD6OjRAqSqJ7swwNv2ORS/2KuyoMZRt7mlDiUg+
tO22Vik2TTjBzxB7Ai6LOXaXWDnYWlri+s6zIhWh8yjrm7JUvgzfXoE89B/wb4Tu5Fk3QGNGbvPv
TA/sUVWgJ6thHMtDPr6+ohIqhsiEJa2Mb/X1uL9+pGRrOGbDKhk77etBw0j1bfm+WK/l3lndi/qw
xiuvPfFE/bYsXTbB32E3jWrp2cjDbBH9GT6UO8WpGGlfV5MGDd4GxIlhW/pb3GYBkvmCC5Q30NuF
i0asZzHw/zDt4jh4nE87mM8B3yLNqP29LvuictgD3PF0bk8BsujGHTcIqXOpKqbqrL+r6dxnNUPP
5TOidD8w0t5eMlfu/UJwwHpH6M7IknaDhrx6HueNVR1aqQaSUSuGijvxT7mN/tdU5+fFlCS5WhZY
gexMcWLJkc+PbIYw0bTi/WGjswwNAoag9SLXgQPut57faX0iAye/YmdX/QDfS6Itiuw9So9y6+kL
Tn6FQej5b68oiQTGB0n85NKTGWLLj4YuuSdZscl+3hq5bGqjUfsstiKXdj5+YBf4Dxb8QoUGgnC/
gBVaP93a/9GkESzW5axkWA4XtsSNXf7WfB5JTHDGJGlGzRqvTmkq/8Kh9Nx2WWmYTW7WJB0Cqk2s
5faC7FQQ1R7G6Ydp/PizBHH3MmiqU6e93ey+f8Iqhkhrhl2C/cv/M9EimPz087IFa4HsT9NJiV6l
ELCSal/dKKPf/gyXKzHc25ba09dGBXspw8f5lHm4VVOBDhkbXvd+e5yCFo6QnE6/woYvXU/59mfL
qfoCCAm81RKj/sagiwN7EVSMV7vmKXUFVclqHZuUBEmmBDvSjjl/BxJOphV7aiMc+icu5OGsoVnc
ndZtU225q5JOBAMytTDIrK820JSrct0NAPB0b+rEDSUXtrF3XXD5VkoLFZPoLFarupsu4oD8LmCC
bJM71HQ8zw8i1q9Ux9QQdsawFsdNnReGc8TDNzAbeXyaNDNiNghN621YmS0HPZ/XRVjVdnBM03GA
JLfjXg++GkAeFbRL/rBy64+j3cFjblJ8Fo0k5cF9BFm0Q3qtHnoY8GRPZEATAkOI157ztyuCFvR5
VxcQ3Eh9/bljWW2tWc+/DmanPsq4t6t/gckoh3bviTto+DY48ljwpRalUTJeydbNE84wZopOoh0C
Q/HRlQBWC4xupPQtHSonm2nUnRtwerXXq7+hDMgy4/mP3OHAJFzunb4bEAn+E6FG1xPuAu/z4EAD
8A+HeWdbQuQCCwGROGJsN3fXwY+S4peqN3K9UOwYBx6EroW6f6UOXbe4DVE/ikaBY576R6+EmmjN
QO6FLFW9jRJT+pjVRneE0dFC5MZTj7NUQ+lLgtI+YfMBBymyxebYvkn997/i5tpoxs8fsB/PjP1h
NuLdrTO5xsJ5mM+SSATEHuLYn7JJEMz1L9lnlR8sWvRYhchT+v9c6mM7qkTZYJ1aBnt9tI/MeU+V
AdjBtoK/Kh1bbd5xIMFnVRYMuq7IGJPxiX5nNDm+lthzXRuvl0Z6RX911KExcdOwVtixqJAmXj59
3TKgKP1eMIxUQLB2vy74DEj9W38wcguz/6U0S/zGPtcLJIgRGvnkxuo8q4DlcxUuPksjANwlzE9j
jId8ohPLExlINghW/ds8noPMS0MK22JqKed+B+pijmhgLXnuKPpBu7NdFGHt9W0Jmv13376mJWax
BE/+Qw3rdqZf1vxKqC4V16uglSdqVqzW8FhhDpjBM/tTrl1w0HRAro+Y/JxnVdwOYI1+B0w3qHXg
jI+c6UwDsYWgOZI9cj1P+b8Opi+rvDnq74UqcNV/KlPMJRUpe13NDSvlT2cCgWC4SotQ7T7N1Q4y
Tb4gkZiifblhhpn5122jA2Bdt5XgO2Mi0QpKOsNE0PvZX/si5PhCYaNWYp9BNb3fItqiipMnpF/+
GU/qPoxIJ+gqmLw3fcW7YD0Vr0M3q5CZA6zmBOZOvFfD6m7AsgwWwvi/gS4B0aRbpTYVEszt3VbK
T84XBG6w+iUvfn4W55rDyhmB1ux+7I3JEY9clQgsjz8XEo0Q/sP9GWG5tYCP2QtIruXVe13WnxtP
BmyP5IZ7tbEsxInv/V2umYs5oz4K0vu7rzC96XUEWl6dGL5fIxyAXn7pJDLOvkJetbv9ky1UcDJh
V3XAC6ATDyqJJ1TMbCR8Ys3cVUwfu65jqmna9ZNnfC6OICVt8XmOoHiaKRBnO2I+/i+XcFSBVSpK
ful/89MRKY7CFfltxQlp/Csmm5RjRk05FF4GyzeXUvqEh5yLtllt9xaE8yd1sWevsVxFl0lW+Eo2
pzmPIYS9to7u2x6TdT8qRzYwXoknaKAr0wFI02QZN27oxet3kFxJBl0F5aGM/rNawy19Vpn5lRvC
56PjEVaQQE6G+SaAFiGivdIbAuGWRG1PMZwI/QfmZKjrnm30UhVa1iJn8pe0u+c2JMf/nBZ53E6C
asiGEHiO2nCyA9VCKJJzomh2pL5Mf2linPEGG8hi+YkcqKPRiaZg51xKp2HWvxRzfofMhtcBtryG
fqdo6lizU/Au2qp404gfLJHrGNUS+/04gKFY91EhlyJpavxb8TtkoeozDC29aAhKHJ8BPdAFjo2i
7ntzsYwVzNLBvOAV/HMGFbZ8HjSf/ltyfoTg6TYlztt3lz8iGE6yi3VsH5SPL5+Fi5FRrE1USSok
5wKl0BOPtKdRaDQnZe9llMYB7009rbajTrTuLhpb6sahqoHvp1uetahsyy0Kc0UyWpQFDk49ioeq
8L/9zChvD6ETePiw9Iwaun1TUdB/uLfD12lzW0rwMm7Gqhm/U847IBAsbZTsWJcCO9oLNT4TpWZH
JB4q9/Fkt9CXm8ck/xYgh6YDWTzwLSBcdmJXDgziCZBdzN9g4c/74cXOS079HVxIFrlIzSkQCTE6
VKnTEHpq30HHLF1j/IJoGHqwxgdrBUzu5WPFUYkuP2MQ+rmSYtksoCP4oXYebuhxAjL4usAmYT0t
MhQr8QEL6LCI1wJcJtMMdcIbgBwZ/5MYU9xd8nYXF5pgeYSfSM/A81ofsFSc7VhLL0f5EurKQqBW
WB9vjgOqN3v/AbUX1xOB6yA7cVOFCcmBzPRB/H+o+QFOJ0qMGdYr6FBGMY8991iuv6lIe/V0+S4q
9oJP4ni98cwK0ItzvhdgVzZqEVLkhxcRb6iukReGRX6Q/zuVgZUqGVed5BbunywNh83P0l0Ceeqa
AWvtHZYVhHYS51Y1Bn0p97HX9lfR+u1pDM00sQRF4EL/OsvNthReGvnXQMnkSoVlLqUQ/Otp0t1a
BBlKGGtvrj80lmctPjp5H6CXL6VH4h1xqMdHZjecpJmcJRhCISJcdQdao8Gz6txKvdtXD0MXVVjy
ezG2MJHXH0c4TuMULpRY6EjssPQCjWNay67orFtDzUgPmBLjUTd17tlM4+9+Nzh8wuq1FORlAnGE
oaWFsVAyuXmmKqT9AIzIDZRlbESKmPZT7soQ8cVmglakatFdZDkDAZtKnzIa2ymONipL48pxJWCQ
X0Eo49l35YF1hIfW6ApLmCFtzDa1NDTz5JibuIHHe93xcjHA4V9+TskZjnUmREax9U0ZtZ+CfvLa
kDtxjcas52Jn/BIhT48QGlXQoT/nH+dRJOxRvXxasLnBiGHbhl1AAI1MlErR9HTeFBtQulTLsOtn
M4tbzmCU9YpfjbHDAk+5DdhYSqawBpAIHUO5febt6muB+xPYyePsqY9zfDujXErImG5iAlxv09xT
Q5kvGHOusZABp7qZ9lhP8elo6eiNO9mTTd0xoPk5pgtcjxKVJgVb2KRbuzgeBTyPhgLbD1q21c3o
aENS2Ww4ohsa8cI1XBr+4H7t6KWRm46XvlcR+X+1fRYhllKnuSl4tME6qN5Iz5vmBHTrN8PAs/Mc
ZfVNxScEaseRWeEUvVttg8TxWlF4rbx6PJaYm8p1l/pNF+1vqXQRnYBnj3YbDoItjYNLRsF9lzEG
7nZ7gc9t9r6BN+31rYlQWCfebXPFtVeXPNvOHE6K5BNggGebjEALer+HkxPOakybSeuKMHP1iYQc
JJvr0/WJeQIDgxZPpnhUk7nE0p58T44jHyS1Us3h2JniDRi4VtoCDviEYhJSiFpLLVS3ekpsZlKr
y1/fOrG5I+NBRvg4H0LXq2fqemCa0SOZ94OjdevNxQz6g0NCNgg1G4Ttn5Rbg+T0EGHvgBlgUaFv
fbbcyf4AfAfYPuvSyVLhcH9CGEcyoz/64701/hbjMl6BsThEgmF95Wmdl0FYqzmgBvg2b9YjncDQ
IH1PQKzDSxNHKn2XnaCzYN7GoqpmUJiDucx6rELRNiugxjkK3ISnB8nPsPY1F9ltUUQiETWtC66o
z2QxSbPAqOL4PETwu99R5emzKz4bQ8J77f/JbWgOy9FPCVS/W432Aads4jVYRT+FRiN5XSOqQ+OH
XYuHXNyVZq5sF3JBipOpOlWTD+GSU1g2sEKeOdbIAIp+BLJPf3um7PBrOB9FYL/M2msBtwVrFGfv
SSMN3h94+I1bAtjMx806NnTc2uJbaURvSyBg4xOWoUWfcMsWsR6qAOBNW5JwEUT96cRgZNcljutw
FBFoWSF4IS4E6XKLiX5f26n7lyRJOSfpOWA5JhPEptSFpBGbDG2cP6YySmm4xhQ2HkZiVZKDtMgD
MePkj/VynCkg8t/oNpYEUw9lNOD9NHTgw5yIIzjv1/fut+dJpT815hNXJ5DZ6OuYlwUyBv6LRl4s
YTJq8M++INmX19JW2LhSykTD6S0z3Yt4m+fb+4yAfWhv+F/+fLQ97rUmRem2pKuvIczuTasuTQgZ
Tm04HI7Ea4nxOHP1jh/mz0ldls7odkmZyWN37cfVen5LoZ2sn49Ic9U7yG+cBkVS1477dcjWMvkA
gAgWBWrQW7DdpCq1gnKQksCAb5rfGJwhsSNsYyUzfwCg42/4xZ+pzpGVR5viCUILqiEIdZ1bZ2t9
zweS4u6geffBtswC4ELOf+8Ya4BfJI7d45bbrEMZjc/E7abnU/+DQ0onHnq1GfHMwDBxUr+WT7ws
zdVjHbMTDlXCA9eN8pD1PrNm3RDkb2qTc+MxDCaGBKBx4RD+q1mygwKNUJICd4mI22KWSrtZBI2e
fRcoogJ5ce8ViFyYQDssgXukS8qIXxVHxlZJHFWoAo6MNReyrOdTqjd48u3fkB6ORVZIc3yGUb3k
iGhjZJ/MaTnC72BHzMSuYBDnwq2ZPtuPo7t4mprMDa7to1/hlGSrt7UXEkxCIfZrFHdoFfaE2fkH
C79W0AukHqL1LK10utiIy0t4p10fIoI3MjEL88b+7ppeCCqViDwqP7d7HerQGanj+nF9C0uVnlOh
3uF0/7OLj37LVLtL/ZIMlDNIkvVI+ZnnYhOGzuVFuiFKv4c+SvysmlFyjPboxcvINjX5iGx5wSzm
Pyf8+7Pa83TD26Jyn16ph0TMsr68JOhrJkaEtUGGPlRsGvNJc/sGGdEbwZxOOlESuD/ldar1K+ae
PFdgwNOQ8+nn0hS4i3sT4hhnAuUVtN5ErFwMsYmHR233WNZwgjHFOqCOn8afg7tYuGW6OG7H8J6E
EVnpb83Bqe+pKjkUsvYMgD1joC2x4GBRB3LZXzi8KcZYupMOQjWIfVoJTmHXhagZkmzlHhPqxLnO
RFDzQTz0urbHHpUf7AcupPnXe25sXiM/FPckSlsGHDtJOG2UDUI3TCjxgWlKXOiKlN2JRUvR4fLa
eavmaj6H0qhduLzRRj6iJKRjB3NEVxni9U1dB5PGCEZCcPNiu1amoMjO9w7DlVyYIAmeXXF8HGRi
LQTmrlBx0w3zCDeFPXKYlpv6o+FCSYue7y5OCoN5SSdLuv3T6vTyu6Td4tEesCg68iLBWXUal7f4
Q8ILc+fXu0D5xvtFdNGNazLgm2SOEyhI3mg7MosQ0xLypUmoEeLY7bBlXs5/2aqyrwsnMwFyO8Qs
nlaAht6dqkTd0hRjlEUUeEronLRcQ33uHMezv+JFPcLNbB/bRp/6xe4RhHfD+972lriy2X7fwNwT
BCh2DyuoEqf3Jalb7dAreYTF4RsB8NnYTxaSJ/bPEMwBz+nEKCYHUxZOmTegHjs/t+Uh1fLhqzVg
BLmibnRIU5P6V+yy/ry2xpI/U/p4ovevSWukeBKIG6PUngC9Q2eEZZt0EOxPmpGxD/efmbLlqCyY
NisnoxEhud8zNSrAAeZsXJymiXm0qlKzP01AEoR25LCEciKJGV8AaD6NvlwmzK/Z6SAtUP++KOmg
P9siyjR+pSR8+dgZZ7PPYeAiO9HeSaAinNZK6FF8/AcAx6ggks/FYWGv936N+e20zPKUwj0qCDjJ
2txRurJFJ68uZf5+IqinlKJhGL1pveToU7aIDVslpjOsklShZOTN/T305kq5THHGzJmh6E3CTSh3
AdcS6nHzoCSEHpbKMam4W8f6GY8oqP5ZqqNwQZztJHcRTf+tnc1VNXt2xQbRd7A6UCWaY4bRFmpT
4PHBrJF5HujwAsmCcJ0bK5juuAIQKdMyAluCMqCFFeNGQPef9EkF/bxcKDxCpYCcGcy0uc9Jl0zR
Y3FBC/kcf5EX7pXphFnHQcxbqWHX5CsxOJtpK06zpuCCUM3+z+MkF9uR0kc3WRAM8GeF69MLSRw5
fmkiipBTFsbB1afTt7vOHVsHP2FkR3reTRPV51lpHeKkxwbbpD9WIjL4uwTUV7JXXzUFF63fT+70
gL1LQsPC9sLJsaGA2Gd0DCxlSK6MDsI0NFiM1xK4yrabvcepYp9nguChy1SeJ67IvQoZYZ03HjWr
5QBQp7IJy6OEZH5AN4DZVPewKKuCQSHPjDHL52jdYnhgZhJffEVf6/bM3/0Go5Y+A1A2ttyLtOTb
gSpDcyB7HvIbIZe+VUIs/jQSsRgwzH6TIlMWb+g6l71BDyNYFxbLhRx602+N27s5nv0CkrlMhORj
vKrm1vlaLXfeJYrdDzTjDOlaZ2p9jhbjtaFIDx/0ecTIdZprp48QQRL3WZdNUFSnLZrc5KR1Ya1j
SckwyfnaAoQKMm0GdpO7efSNo7eGENbouSAAN94R8/gfcwbo9qDRl/Cx3X08I7SaJEGarmsZsF3p
4OEkqmVPK4VqicIItXsdk5RsJTsH9ZcbDS0raLgR8Mowuh21VtjnfHXq0KEhhgxHU5XIhKL0zCxJ
bRdcgDBwOcDo6xsvEPR6Y3kmsUChCYhDOts23Re0Gd0No82gSwmzqTwc9Zi6p+2Dtq/U/wNzFaiZ
gLetdoD340pD2W4Vc6d9jbEoqkwzkjTkaA3XCGL8sbVz+wFgjx5d+oXIoTp/xA6sNvBykLvONF8y
Dyy3py2qWLsc6r8opIvXCtKeb7r3D4J2bwliRbu1c+TU7RzWYYlWzgJbd6WBCl6sm9wwXlngPt/H
ix8y1QLYcs4rAWM0GAdLnXdd8MZgDqp0rfCbfW6CH+qbv7njVRbabj2hTKEq3KqoJBzW6jGXp6+S
DhtyrxmMfbR5d7tg4IzUZ24oR6xwavnOo3LCQ/WmHR/aF8Ghl7vdpsVXiONIIx14XUU6hmbwX3Ic
sKJBdfjIBNrumzl4XSvnbh06dUKFq2KUhqTqvGSoyKEITa4QXMaZfiQgrsWSG8Qob9kNMgnJm+c2
f0har82NcCtNVGHR7vaznCUHOSLr47J08MQrqaiasNJAito+V56SMbgMdHkzxLEZ4avqkPYjI/Mh
omZ4wgKFFRZMhpNHRJw8VCPvwGUyIZfSSPvnWk6BbPM5EpcSXOD9qsPEL7WvBFH5rg9rjKio8r/3
n7VGs6g7WdIRKXtOYRFtwk4r64T1fk2Y60/JocMtxceLEDoVlQTVaotQ/JzZ0oI8YGQX0raRcgmm
Dx41xJeuKjV6Qa9Iek8wYApYiebw1GmbH2eD6NkbGBNsia8tKdPG7J7OohTuLUenE9p3IRKADqoc
ynuvXrfFrg+H9HDhP348xN8zjUU+QLQhYCz7/yDgCckGhJM9IHmZBosMjMjIPpVKnPUITDAeDOPs
m4VNNGRl8urhcRYHle0qXX3bQ375Wq5h6kAwcnEFYS6oMDU4hJkeW+umrBgMIRg9K70u3yrbFjwB
PSBlR/EKXCq+DtRrfrLMSyYn1dCQg7G9dcn1hWcq4yYrqCI1bxZccntEhIxeDODGUG3f44vFnhYw
nNyOTaBPoFg0NOrG6B/vp8HjYz93Tib9EjEfC6Fk9RE+ead2wpo58sN1LxbTfrBYeeTneQptGFrU
50JEC3SXIr0XjO/TTemObautXrSF+FtFMokAYNKUb++oF36pDZgO1+9aI+3fD6uB6OR/TOj3/DbL
V1F2AbU4MvJpCJRN54EhNxIcIRVmreSdxWiI86GKn1yPGEyMeSNZfTtFLy8SM5AgSJLxcw805tBR
H7MXzk3AeTAXaDvKIAHCHQ6ova9cCbBT7Ab3chocMbIRPu0B2lDeTFIdQ4VVU+lwUxI9HggS811c
IVI/wbTwgTQv/WemmYoyCvw9pFUM7lgORreweCaF/6nNB6vqhTo52K/bEhecHSBjXMdhrUok33wv
nn+UZc6FwYu/TekuedhrawJOVC3W57zQuUa9e5xwD9U65wBccWd1NgePon/BIf2q6yF6uNRZsiFD
aQJiDPIsx67BcvkgO0a16VHbm2hZpEkLS3j5yOqKTpt3mrI2J2msF3Wb2sLH2TjN2hsJt2C2q7/O
g+ohPZ8+XkjzGR4birFpqeiY1AUoXusRHTs5P7SM2DWRY8KOXgt2UL04pZaE3rTHu+s9KHNlXfSD
Bnj+0UIs+HrUq/dQlui1adzxq24bGHA64IKxPR+xLlHJkCEABAGxduLZhV7GahzHhBRhfJkfesWK
up5p64xHzxU4P4tUF/kFRiq3D2VmvSWWQZ7Iy7I6exFVVa7d7NV+zm4aMmARk1C/pwnqyifm1O5+
qBUF7EKW//b0in/9Lb7lhdsp/IZpWWAxSlPSOH9apmBcQMQPWDIL8CXtyU4A2N0JNw8j3fca2dQS
3x16RUnQJS5OyG0C3OvQIRwMgudB5GVO8QtkuYQjP4byH1AZJEMnPphlYOjd471vYFp1v69optrq
4PPFgWUF9d5ZJIM4RwhrN/8trhuwEnqm26qlNgDZEyDoXPNiRRzzdH0/iDGIVzdtHRqLPdMaz3+8
Y4jAnZI9djKSbZV+dS0wm+dZuqqUn3JMJJwc1cUXdOFNJM/OHFeJe29k0JX1YYvhNtFtf6m+IXHM
PIO+hhRVhzi69++7TkQw8QgjTPDHSdv/3bgF8MUFRW1c671B55sV4G3vmoMaA0fpI54v72LC5eZr
k10w1iVBUWb2BxYX5HpWuH5WqiMYg12VZggGvaDuSQqV+kYVNULO15675uS+7eFpXm9p7s+e3UaX
XsGrjN3q4PS4aI3BzWJ3QNdRqpr0cAUQEXbPbfRhu7BmAm5g0TbJi5VCjYzGWk26VFFiUKWpErr0
D1y5/Og44SYs1XFB09VAhETi2bGsesL+XmVzRfr5u4nxMs8ozlnQinJGs1obo7mAsJhrgzVbK3vO
RrB6cU2rEkwpr5yA5IbxO6u5U9RhgeB/N9nCrULe8B/0lKcLZwtl8G3Cf8OQe0Bfi4yskgDi7Ld8
0S3kqnXS7+3aUHdn7AuZmiFxOCpamMturHWQ1e7UEN6MEHBiDC5/RTxAoetXf7nzJktFQI57PKr+
wMWJOFID4RV+1FTUbgMoJXGTFVe4xKh6G7uL/e2hT+1jYBC1lMieRRNruY5CWe9ghUa4OOTTVh4h
3ywr3MBV7Ev+ORVgVu7ulkVaN9mSZhYUmpDYCI0pkOjzyoHvzI07J9PMwzYDO7oZ1KzE7YFEpqAO
i4TaqFfGElkPWOQcr8CUCZY8nte5Bm3Q/Wj1s4eosgH0kGYS63zinA/H5wOjHK9BhteXWdwjd0Lf
cve+lu5KUv69Ra1XeOX76PbLHmKJ8cyjzAG3wHE/dDn02b7BwxF1p+lh/Eg93Bo+FEHUar5AUhY3
4MwfftR8jbZp9CGnREk3wgONtH4FjYTnkrOPSp4WA2BTlbhRyRwfXy0I8H9ryuRzqTvWom91jaK0
hCyd0bNChFnmZfowSteRP+4YkbE/swHZqV6C3MLl8eDmDvEZusYBZUt3S5f2EWy82fHY/+9OXG2t
HUjse3vIIINnl7deWIArvz0cWOAQu/LgYk1S15nKko4WggSNnBkAG9IlG8KEch5tD047jGhELaVh
1MwIbyxaVg3ZPPQzrpbs0AV6crFUyKtCs1krgcQ8rx+kILdj0X2UVmE0W6nwfcBox5ri2gCvwIsS
KaWf6vUlP36GjRywBKrSyryNaQkfoxQNgGFDJfP2yYgfxZSkkp9GOkAwr+Qy/0IS9a4vzRYqNtlc
cOplo/CabyEgP//nuE3cNpInVUn99JKFs65zCkytz/36wVFCY0nlfN6bZ6zEFZUi8XJsliNF/dfi
TFvzFgwwMyOUjpQ9yUNqB9NKGmJpAm9DGbEtgNxfmrKQ2enspBP8OO99cqPyG2bWfg8lL7Uy6xDu
a829w4B53dHBzk3D0k+Fgn+z3jS1RwhhemYxjquf6/kwRgVyXA/miIZR2jn/g0ZcGU6HRTY/G38i
8rKSF4FAQZ+6O/dyrHsA4fdlO/9kGZRekRY1RKYtok/lx4l+AZYPu8iTGO77o1Fw43tgkQfuRbKP
0eFLRz2ITG/06C5pUDDpinTRJZp1bD0oUbqWpbLd7GaJMP3CnD/By4R/eIax77Nygrw1QvLsUiYg
9Yw9ypotP52c/XGklY4zrzItelQbnPABJY7hFjDieUKhBoAVMQj/d8WL2tJKz2qSCqgyUx7t/f39
qrIlEcf2EPifhlMOAGi8WG6e96kuid/PBScxN8rtvfR3w8t/WNfcaG65Kny1vpGcZPHaY3ltnDXN
ZW/1fp93viIrG4VKGrUiOL0tRIpaqHun7CfZ7vRpTX4/Eq47Hkg5RTby8n69MyRLcud/TbNG3nKy
wrN3w/6vq7T+ojcvItUdc6Lj40Pk8c7/9RWd/t4bSbn1yt0NYDZKYhRuijxT09PcuqLTRuDMvBDF
cayyIHjYZnjih7d/cNZSjZMh+wq2RAuj8YrONPHwezrLCofTAd011zlMbty2ToVuMOFRVZgrrWt6
aVywi0JBgSbeyufqx+6rx/OtpdnCExC62WVj/90Z+z5ZxHrlY0koUxUZgJ77aJD4HZ/L0NoV8gdc
Tqp3vN3ZN+UZeB/TgJFXTI0cqksj4ExaH9DMKvDdqt5VvHCLbBltrS/SsGq/Sg/Q6Nw6g4THdXph
mKIBwr7iEBmRSSq9OS7EqZbAVEMEJ1U/8lIIxnmZjiMvsN8L86433nccM9HTqaSBOeNxfIMi++Bk
ON9kX1dlNq2D6Z3/aBaMG3MSEjF/MaEMMRKnVvLddfyETKp3tRF2Qr99NrgjJ8iY23WmHWUmWBJg
ys+9wX0ffPM5IN2jU1vyUQ3NsHlrRdL0Ufu9FjghkppMf7JyNQoHdxGyfM6amITVHGULzFJpaMjd
oQl23AJIQvG+ircQvPTAlTHhIP1arjVkthkkbPakOurtfqy/YXY+Y38RNkAtAkDtiZnESAuWVxXN
VCZM3GzsEE1Ax2F12EDoPYFG/OtwHBukgCrgduj5AElHPYIgxeLnZCgwn71o+3dTD7zowVS/6RTS
CYWufXwEOayxGt65+w+cb2dhGb//RccrIB4Kf22p1B6dcgDL3WERWOW3T0UnblkrLolrbgMnBYSG
f65pxAZLCzago9duXzv5G9IgDsx9Qe/QBJZrRx9bUxVKaERtFfC6Hws6bKLIe6r9yKQRwIB84dxD
rb5tZ7XdfqYSoL2LqJFFrHU0oBGhQAu++/sBLHcqd7FzEKFOj+UQVyJPazs905WOSOK2gKN+fvfQ
L0es6kv1jaLcOaeSymrgtZ3A9aBu20pRysiFRzxxKZz//Lj8DQLX77wETP3faxgr4jyrsqTRMUUU
x19QuF54ZraPV0nlBUDOBl16IntTjbtL9amQJPflNaXVP9N5vmDKzt+uimRihzush9Y60wf+loJL
JkXjZhL1+ZAgORGTbDLJck9VgAYCYIGgGIkk64P5E+ruQMZpgpZaPJMQsscdG5eGva8poFe4WtVX
rl0cz3xmrrxEVHLZsc4L7UT6JUxRiB/ow993s4QVLvOjf72tcrZQK82WqYNBPpdAHiqMlqdNLkwE
B31wvOkbNvjqQdaRoMeCEAZx9C+94JY1hmc5+BNXmkECyHYpKt/xy+fTkEa0kSieIbOiyP6pwBTi
+ASC/CENV653AI+XjPtIaMlNgWHWLXCJ//z5fr/TwLeH28s7Pvbecdnu8nhge5MaRNm66Ztz+uNq
tJehiog10hGZNhKeUu0kP0g7+7/XDA/I+SHhEHn1nSTRTkC95RZIQqDRnBUjYCC3LRAfjgTfMakw
OHdHFNW4r7d0AoDWApOaqa8HOaMXA/jHgpGq1AnssktJXen61nDF1MQpkUgbHTvUT3HXbHfVADaN
DsbxqLTXibHeXLNYBPa3Xfl0HBB/AOk8XAkNCliHgJALndCTGHW5+Ia94H6g6yqClEN1oLxQ9ShY
4tZD82Y1M4SMSklVtHYosFWsqETDXOPPSY9RAbRZZLWRNeaCrlUkj+FDwgJ4I6J8e+C5HbMsKfZp
0nDLPLkWpS5/uoQW71LUNVAzCkFJiUWDi+Xi3ihAI2Rb+Xzy+IRaJSmhfPPWRLMq2QFyevBHnk+M
Q/c7/feddqbCqxQ88kd/CjDlJIKGV4X90UzAlrXy0kRA99aXHQddP3iO8vUOgq6VkJD4Y4gTAvsA
ccx0f28a3wuBQdLwHBLZiISHf/5+weOHijFTDmgmOF98RSRFfuy8on/Q8YVPdHwMgPXg8rXY82YJ
fxfDJXte+nOvZyj/8IowNi4Wk13M/1XChvSctOi8WRuYI13OR4x9VcZ1mkF/buWURJCVflS1fIkr
xtUXdH7dhJn6Ca8EuW2w2RgifBlx+8uZyecINe8N3SglNBUSIWCDFLVkLpTukY1ug8s6YkDpdOGB
pLuIdQFPMH3i/BEy4jarAHY0SjoiclXRccz8mj+TC/DJNRKqUBirXD9ukvMV/TGtm73Tj0sV9On2
Z+IxViCnoDhAWbujLUyGsnLC+Y/mayxumqJnpkXXaUWkaaSIu44CHrR/6ZkBO0IP5zRCzV3xkOcu
PH7ee3LxbGa9RSXOLga3oj4GOP7Nzcc2EQVzOsyU0OvmoqiJzmEzw0UatKauw19RWimyMD/p6JqA
raidO7QSWNDTRPrmj/RlcIYech+hgH1oDJiQG7NhICvlfaKI+7MZlw1FUOvc0NC5fonAjkMjm7kR
Dha2kjRuz9vtDfPgqkN00yPx35CZe4caox3orPcm1HCphv+c1j45PyL5HAmwXkazzb5RXggcKEON
Ombd3DiVqdZnTW3YlpEE46NEGlb4DVxP1pE7gyuD+nPTXb7n35iSgFsk3MqhmcuEtZ+DD6jxo1wD
HIRho+fqHg2LGXnvptwJc3bOxGaNQLpHewGqn85d/Tpgb9HKxOKkQ9OkSeVhA1Ng/QuEP6ZehNTf
3ZO37JWcWj6MB6Dl/7wKnykLmZvliCvS0jgNIgk2sY0+m4UN16oIlsWZ62dwwvGIFW1lmrCCZqSG
2PXbtMKzLf+duD3Uw5jJSMP5niv4ats57IAYaLvQ5HxisrnP4oJ8IRrTlQU2q42+tUqfVFpfGlOR
D8YpWhtB2AXVdDx7fMD2e8YjK++fbkGnv+/hBdQ5L4P42um2h3g2iX7IeDHLjKQaRqcH9w/5YwLN
Qqi70jye2QjxfZze2ED23S/319oSOIgcqX/o0+bUrB/PgXsEbyBXfFGvLDyHAxVPYMxIH30wae4t
UDSwIhaibb+5wXZhl7naNONQxazqLLU+IRrOdavzfXSXfTN7wUdFmG2cGrWhvBzXQ5mZs5VxBmx4
/9eHMWsJXsgxImeXXABJeArNYqRgF7DKpBuBjof6uggXxu8VMaZsRN6Lp6dyBGyVnl1/duOSSnZW
R425Sn91uPCDTFmfqAgMDoTXtKl4KIlaNVCtAwqbjHEFyt7O74AaF2alU9gn5EYA+cqI0pJ8UuSr
37npBp+VdFs64lwqkd+pZXg8Sjozr3PiZ0369rqxst8DAWh2kQmYFUXYz+QQ/Nrbhvuw3MSkRB3w
ONgXk1EWZ90AZIGZ8mBE5xz0SJ2qZLedSydx8XLHcn8kPlGqvrlwoUnTwz3G+PXAK2kctbHTh4vX
yI05S7CLB9OQjcHgqcIxqh9yeQiViF6WSzA+nXNvosn58i1QZeYr8F24PpdWhCFULy84N1aABc5O
R/qiYF9vQXMy3Bse6vmx6QRx/Z9hBGxpUN+ejlR2KPfPxBkGC26EAHvrzHYWKgdvkOKb441fnY9g
9OUXHeO34PGHq2bm/Gh/lEt9s3EEcQYAFEj08cI8yp6X8jipCu+RD7c2xEr8AdCiTycLsJRCttBm
kbW1fwB1xv2sdK3mCSKSyANm7gIWSUG1j8AY9coaBecZmmszRX9fqdZzJUT83VGMRcs520b1WRAe
u3L3YxBexY32SqG0PBKvCBTxLnZqQqlYULO5fMLm1KXdoZ+fAuI2fhFe6fAKfgodLJbPkuar+/pM
4N0KSFhBae3XFw12rssvaVN1jNNuCNswB5hdoG5HuTUEhyxQtU/IwVfYHlqlu19W8Ag4naDgkNZV
lBbyigbT8z7Jx8jEJPvC3oI8Z9LneZzUg7EtOltl+65J8SXYhS2gDzgUGYXsl9IEkv1X5921jMsL
LI0zGmdfa/pl6OYPAyoEfr3/kIIjbY6aS2jkVsWFJDSEBZUkOxCUXK+zydLr+uxYhyLF9liOOg7I
eJYPSUPHVsoctTjWcvapTyeCHR526UMO0fhkFAfdhYmuUwIvM9Je0YaTijSBNaRvR0jn0I/075T4
w1T+4Z/KI7xDYg5WDcIxk81/cY/FmVge9STpC28kKqc0mHLLrr8wXA9i1Rx7pKcw0SIT2KOhGW0U
B2q7kBhWtwM56WwYQVeT879p5hlqTzn+6AovE0Dp89N+rnrU82HAiE+PhUDAJqrs6D+Elrn8QM3E
qVf4Ft/EnsdE6Y9AGHoaajTBhpdOp1LiaiD113kPbcs4x7pzAcPo51oJ/StONKB/NRrs2L0qtrSo
jr2Evh/OQohek03uZ1c61qrlWj0uvuhsB60HmkG2LQA9CzbklUreWPMh1xu3eJYZtZzyiAPZlz74
u1RD05rmWtHeRE/KvIfwqHJ91IpADWY/R8xCseCVjqvYjdPvR4a9myNUwDcUJ6g6uIsI2OW/4QMk
mOmEMPJ3ZhbsgER0zhDGEj5yuq5GJZ7P3Cw/1SBM0SDdBUh+/EyFe2A35WuhSzVMXOMZEiiyz2CQ
6MxCIAEMBfIg7LYhDcVPqSb3GPzls3Zuc0qBL02BMtW4woGk0S/7uyFUjytfUXkcyhyPvUZxllGh
u2fctov1KTmUOxyWnmwwhWH+3G/nH1PUKxc2/0aTOKSy4CGmbm0LRAPg/L5vkJPqHjYKzNit30C7
klQ7s1Fcf6rfFHkaQnkexIEM8RIell/2tOe3ukDf2Xx/Md/XYOaDVQflWm4wjBs1IzMapuf96c5w
ttI3h0rv9AsPqyA0yb+g1ZrCarXFL0GWlKNxOJ6Us1RNu5WfJFpWyCWheVAnCEKthd7UKIoGSg4T
JxfXvxur2oe6YYCILFEKWbFXn/pflMf3zhZCDqx0vTIOAVC3rkM8+MhsMiHwAgFpSkIw99GQVXdB
ZApgkPkM9OgJru5nppqpJe6enCDoG8pCU0P4aRJpuo5wW4TerHdhH2cb5RQq7KZ/SQCY1/3Orr/8
D1SfH375wgKYHvaTJSTp+fj6o+X2fyDIH7bEBHZEp/6DRkY5vmENhqzWGoRi0GVuFryqWKa3rjxK
Bg5pAQRJ2Zdsn15C//7RWVsdA+9piZ49N3KUjVi5krvJ+oWZ3nWT1uKri6bponp2mp7enDPN2Gt0
myAFOnAD4iIO74MsQQFDam7///9LWc9QF5QHcnLT6lhKMHTd1/e6EjOp6STU/tBQIfPdftT3bmWP
OfiAM3uitucMavTHNbSg0gILXiCNldP1PoBr+zSIbGkAarremU6k28OklfkubD81do+dKjnAkuI7
+OIoiJEyM8nbISoQRgpphRCepPUx/ro7YvAQy4/8ZY6w1pInPRsFgjGJ1EawKEFeLV9nPZe5p/sI
5z+OhGKA55n8DnSaEhw9buLTy0cphi4IfYkrp5o931wqJ2BAmpu8FJsJz4igG4IzJuNW0EOOiQDQ
CA0WbaSqFGjfsqA5EKIpFQpK4FS5PqG/6FOWGawAFlIJlaCGbSSCYTEwwD7c6lka9EKvG4xn3BNX
3S5xixNzC2dPUcquulorMvwEYF2aNjyfFtIBDwAM8gyo5XE1rk6tg+vomY41bw4VYCMdgC1gdS2F
xPv+kd6ZvQGXnjfxC0SLfW399DdpfI66LtCMh5Snlz7QlBVT0otKhP8TWHZ4dQNFCnJNPFX1sGf3
AeJfhWRYIQZquX0SJLTyMbtAUD9g1xT5KBQVjhoSBjgffdJFjZNAFI1jLio3D40eK+nLfRYEtPr3
786g3QMLZmBTKVfsEubH9cRFjW21Li+WiDQGXJGeVPzh3EutbVX5AWi777WiNq0ugyoFd4h9RnK4
qKasoJS4Lu973kWbERADKu7ngKXbkl9eq1fGAPWUxjxI3oJPzxbb4R2kBNF6oUAEETWvUXs7WGe+
Esb+X2R3KM9LG1P3tTTwo8q2Sir0lyBbO1UgubI8SngvdeApDCVWhOUL/5HFljw65p12zmS9Bmq2
0mIdRJrklQxX9joPFgWET7iIzKQBagmRG48zBST7h9kf+JtYkHQPb8F1DJ5wQ/9s/txu878plGQx
WhgSuoRA0l9KDvvosljNCptq+LjNiIhZFbG2TLxIVLlUwbnWfOHga0IFLiTP0QWlS3jiAOIMiQ+F
cpBKu6YYCcVrXCIe9aK9u3zDr/bj/UMdlYtYfuHbm1q25OnuSL/tSUNgTJNnuhBd9WSroE/z+mId
2jfG2p/7jh6blu+AVWta03pu9aR7CSBgrdbHMIQzkacfz6jOFOEhZoaWWXHyRe0IUXuvBsjp1VE4
/FAn0mLLdQnDGguPF3JAhINzgewTsUi613F+9ZZqrbF5YAn0lmKfEtfPIrlAxlYxwJlxGcQ6en/t
YzcaYtH+ogOM3qhlLI11aiu+lnSQmcRWlb/hA9TkCebFTWxzFo6OSe0/IlHjnrbxJnI1827KrOu3
84voJqVrz+9/xWJ5ow5COrNGUywgnI3N/ikhyYrEZ8JvsJfpFbEnCd76ucRkoBHOuS2z9m5siVRQ
CZXEkRVMPiS37VzdFudFD1O77pSRAz2caCWHiELxBX02gyLg+3NBqScegVAAjm56FgVvSIQkkWi1
Jh++71qVb3WV0reay/mCh5eXat1t5p+48aHZgoQ5/YOxIS8AbQGRf6p2bZ0tCheBWtw8Hxac3KyY
iGu4wN+eP3tgUzpeoqw1tHpRadAkCcS8eJjirPVqrD4MHpy8CvExGkvpo1QPSELfT2Kjb310aytS
5jHq4azm3lBdyRWfSeancwCjacKrkh1nM9/I4ZEIsSwywkfTEDfAxFRFO7+TAv9gXeQsCrWo0vX7
fTXoyPBGzI4Xe7swEIgyBJD0Rf/J0ags9xqHXL9rjzNTaBLjaBJFkksIMkTV0X+OtIhaOHHZEck8
cw+BlCzYROAHqDMZfQIDcHQQhOEmgXSL94eYBQL7icXDX6OYJIObnPDsSyGvjNYygM9NtX2xI1z5
DBE8Z77Z6DGE13fO8HCn8sNwe3/fkAQQ2lKHEMhoCMkJBaBhQkuGGZM/n5v68b1sfe/2XqPPMUnY
kAzKpgGFXy2ADfBeLf73Seyxr/slg6yzyDP7JMfXAC/sQigunZOkbncCmylbEKPs5rwOFYFGTsHD
D3hJfMpFZhX95D4IoPVtZ6box2UCrFZoRRBbmCVo5gN9poE9YqboUJI7Jy1O6dN4EF5ap9Os9qkI
zlT6iP3ybIvFCecbVxFVLNMp1ucMMhIswOhRIbeWbSqA8YnSJv9hvspOJTyjkou1YI3+3y7LemL2
T1kvdh4FsVMm5pxES9PnT4yT1TPqIj0D4CRf9KqfMyrzyGodesxZU+6etbuQWGDH1AV9EMvlvje0
rvjrbMcuLjMmIp45DL9qL3wesnJkhtHHz4d/Q2UTKdSxn1Qe/XvKe7Clk+wkd4MH4TS5EdXI6MBL
gWPJK6dxBXXHzzmfYGWACnCQItNr4HMXZ6iBGHIZ6KXtlN8KnXe0DXyA6nwf598UrTRAsE8WhnRT
V/W8MPse1FdktzZD2/iT4Jr2g3f7wkT3043cWomSTPf05F3huzDgMKxS8dGa1OROL6HkfORyYKKe
RCcreNZXN31sM/F/3B+ax0J3RCv1qYRHrB8P5l+lOQQgAc4ItVVEoFNaIgTxN9htZIeTSWeUdnz/
Y/36vM2GKbih5iRdgJJs5t5+z3vMcEGIovENM3+tOBxB9i42Pfbq0HgcKG6uxV6Ea/wPX6CLj34y
Xg9vPNjypjOsJqECZSwz5p9MornyKO+AOSbHBRPu50BVeTIHuVsvoRzOD6g9GHiyaPdrGTDyXAli
J4vsc6bSl0UYQv+Ide5jBkQpJ9oMGulxpxFrwkQsDvWd6dcG3qnRX8MHQD8QP0GfJfwVcCXWsnCo
wShv95QRkxczdIxoLy4wgE2JEtt3qgQAjuqeL3uKAnEMT/phE347jHpE6BMXPVHPNBDEdy5hXucR
jDFda7s2ju7fzKGNWZORgZe5dpDydtB7EsfCYyWstaodpJMtWluyRWYWSAw9HBwEJJzMKHGHPsqj
t4WMD3OosiBlCSz/myY26daZpk0KS4wsFKNzxbDornSLdE97Nsm0qkDONDCyIm4TMF8AVQaTApYN
FnNaVefnm6D6Tphh/9np5JmZ0Zhaa9HQDkasMmnw4L09kxyQCIAk6C4ewpmBDE4aRbUrjODPHj+n
84BsXPKbyR1d2mjFvJJVA5Akm9Mj+aXind+Z9w+00KJfbI9dvYjlNoIl8oZw7dEktQ+bxO0a33aM
j6s3hgoaNP/zb76bFlbVdkv9q+zNeHxeLoJdWqeNsBwVYu3GTATnyR/kLDqxDvs/uj1pJ30eLcgb
M5Kfyl4OjPh2NQ369RPTdoltnfCR5mLW57+9Z/aYm0I7n+wBwviQ7gG82czluCn5csjTlpBYtocU
YgYun/jIlca9eiDN6GmifLI3yLu4hjBYBrhbSUepdG+D6e8u/BGb9I4lYaRM7dMNIBmuEOzvaSeX
2NzYD+QSSA3YuUBlBZTKFSOMsjp/J24M78MMUv1+VTz8mAz9Bjf+vmf7tJGBtqZS4ysSMCn4Sc3z
vxwLBQBxYUVKeZN8N5YaPQ2fmjnVwMtT2e4TadNQstzH7lSq9Hza3mJbAjd2ir4hOnDmvDTi8MCK
3VlV9kbINK073EEGL2hBhjXPd64RGh4UK53795SHttM90p9ss93aK4AbGhWGctz4QPPpmKa3HS5H
XGCvUqOTKoy7qN3P6KTNXsvmeoLH4XC4UTOmrDr2IZfcIkTzDHUtaQuBCkOfeeXlNqDeZ9RVRb3D
JdYEUGJ+RQpmtNd6VvecyzLh1fc2lC3drVzTsPT17JxdvhYPU+M+0/QmA2BZBLffhT4/VhmdkxV/
tRoh0i4SUe/TcTt8T+TIT8Fj7AZvnQdoYnF0TbkNPCg9aqRAUL7wfnP8SmDHBgBAnv11i99U9E9T
u0SxKiJNAxstR3nHFfckbQqzMq0a6WrdIEiRTddm+TG3j+m59KGUg6WAtHMHG+fs9SQUjtVfo7Oi
ZqQFAr+yKpKMYbVQrDu6n91AKdANGDJjKbrjwD4SjkAHu9vGyVcJ6amR072ihwaynE2pFReaF8hp
2wzrCt4JoI0aUDo9Y6PTyWN1K7f8wIPWyp3eR3Qrg+RwgK0BTGgFg5spVecFgSb3kC2bCrJaXXU3
BZgJU8DtNFvT7CS5fdizW38YUgWEFPYl/wohrHQB22HjNxltVaDtTAQDvq0lQE74g893i3OvYVkg
VNCxn2lJMJg1/TzGhNPxXpWL3o2xpvK4WPGyzP/oziXbIHV/s73m0eBWAtgbmO6a/vs2OEo4eNN0
LOfcHyOp7/syCVoBpS+TnlLKuswRfhJAUXO8EmnKfzkZN/kT/2xu7HdtbdGN6pxsYGgwQBWnwKmF
opLN6e72Xv0Y4KQZ5yXN2eAi9Vu5+S26awJRvk32w4m8i2MY07+CgRYeOrhvmD08kBjyE1rX2O5B
gTWRZnpf+Ojb5IPx9HWIu1UeR0qS00rouhQhYumYEKGZ4Q9Y26BCUHV0xnwnp18nB4ypj2rL4BQp
r31r1Fpt03oqGAHvG182nnIVjammIJhHUErSEN0hENiJXEuAlwyN5MUo0cZPB2290wuvXQlayxGx
sKTgCYKakdtHgpCK+Z9PQeNcDuANzfd3RvLX4CD4ZIJqJfRxCsOHNPbeGbNdQkcpeiebVi1GqWCv
yhebeHX2HxDEe03fntMrxZUDz7yY8imkitZPqtjyPQmhdvIciO8JfLD+TPcYG19sCIFu5BIG2cvi
TiZlYHgNtYD/2D0Snimav4yIkzOw3E5rmbDnw31N1p73UQWJDC0M5PTYQqgHxnE8OwJTXegYQxiq
rVqm7vFCJSqmmzITRqfwiDO3tsxttrIup6JuaOjQBjKgSpGtrjrJc1Glk5bLF3EPK1sAH8tCZtL9
myXXyMaxp/oPqACAuyV6KZ5EljZVVloPY2G5VTEVlHKynxI3egCTK0drB6QRcwNjvOu/Jud4Xxv9
cvzLolaIcBaU1MTW4/X64j/TgpQ8SYVMtaqxN3jdux6I4197fR9fYXdf7832EW4IlnzmALP7PFA9
7ujr8QdskwVmaDNLEHG9aq/j/RSar3xVyVk1iCFcOKGINIoR01k9vjYf4Igtzoznj72/mFPtlEkT
TGoAE3O4KVHdejkaxsDswERz3YLpCW92wp8T0/KdU12F84xpIrHQUMcNj2etZBML/yTER0JpqFiC
sFT/4+9pcK/z+tGYVH7ue5tV6/GWY7XXSecOvutGVNB7HJsy4itXMjbadyjqLwC8KXVgcD41kPhz
0GQrfEKDf/AxYhfKOnC18SzjsctX8ClIzabzdzhLOxijPMWFnshRxCRFpafgShD5og4myGTkY6mD
g9tt07G8IKUAMcWl0T6SCpmnX2/qKzPppn88cYlBsl7Y74GuwSLyXkcMYcyj6KG95hv7xTXczRq/
acvrzvOA2MKPZ6Y1Z5580F0wal4vItVlPfNI3vxrjCWZuNSbIRI4U6SfXW+J3YDZa/yaZRz2Cru5
rznhkvkiauc9kQlzmbHs4lto5kYLBYLci1jiQxPUiuUlO2JQjRzk0Xy5pbCiPNd7dd594NylGfHo
lLFhgDKRhEB5FqqRLHPnG+H5X6jE5pWgs88o2awM1d/7g7/jf+RYtmqeYLDo+GIc+mYhVK2wr8L+
+XruOuGFGVqTL4njBa0FjvFfYUXodi+qFFzhySOE+FDWv0Dao5+IXkoSZFuHCP72ALtxe844UoKE
GaO5oVJsad8ruFwsZ9jIe7UUMsfRh2UM60JjEy+KNjXOqz4uaRZTgPhhvHtwuWQ0buDae4nfB5jM
GpSi5spiOFAbtj3PBZJouJvso/8sfKp5WUyHqcfATfmxIsa25wDmEDuGvVVcnCkU/WGFwgiEG41h
rf9gOyEO/vuOj00fPFBhiyIEzlZm1n0JBzrDRgZmw7nEujusW4Ofj9VP+zNyjDRPA80mA786QdEp
05feNrUreCpfvV/diaNzPH+NJEa6xq1Fsntc8M5/qFN+fphQo2GV+UKKGjXK2OLXhbVkE6epZTtd
rtF2kjiK5g8WaphSRysXRpYOj8h2QiO6BaOMNtssGdLxvwhqewFSFglNL6OaTUbsp2Ka2ZuVrdZi
95Scy44zN0VfYzKDAcMgTKLN8J0cEd61pCLn/s7FLLI/x3Rbx0m7YqV9P2dCFmMUXe1xn/1f+QNF
wPcINWta3e+YzA0OxQMh9UIILHO1sFnFGZgMb8eyvu3qg2edAmoV54uA3Vro6u4jO50q+3XqK21m
9Xj2vuAEaaRuVhlh16HxGv9QTKy9TTzY6fNExsDKulJijbFUw9rV0a4pW5AGTcPUelHQq1DlPQQj
fwDdb5d77CZUrYEFNwA79tzftYCnddb2GrMrKdDVsxQUNOZ58HWqrzfGX6QL54NN9ANkTgi5jhhs
CnlASQnNoQ3zCRcWA9ZQcTNfqSKdo1kkBkgHuXl0U4CGXfl91UdfNlxc10hG/xSIPJUb6HYthu2e
1iWoqDO2ENCAgsovUPcFHvUm6aBKW9ZkowTt6xmALlZD34gqtT6pg9tQQ1DD5Zh2MF7Jq9oAyY0J
Len24zgvUIY03XfEHEgGYUeySUwPHrHD1qEomvPAAFSPN/1T1dzumqQZajWt/Sd8Y9SbNw4aSKmG
sA7Ew8Z6sGjUdRWvzVNP2JZLrTtHcnkecDzRdFA9x1GIZwjoGfLbxwzflMeY9yCD5U/3w7Ie4LPo
Do7GoWydz2cyKvEHThwQr3nlERjoX2BxryFtYoaqmO4T57uqMkqPuurfuuzihiMOYzWjWB4Usrf3
u1Kisyk0zZGBzRETnYG1p2iBmglcVcf20qvkNYKZrhNbWspDDjE8oOgkLcaUp3AdWxdboQvhudrq
NSw+07Y7QfxJD5wFvhtNKLr1lfGYH6+CTcEyIFNa/BIsBUDbt7yBp8xezAKKTHsyHiuJ4CL/Kz48
a/irUwS0pCA3T6dZTspcoebledSka7rJSdFeMlDb35rfvXETdi/98RGdkfsSFaSNm82DX6yzYHys
tRoUDhW6OwEd9zSS7izPw8Wnz7BocTwMzMV/bnY/Vl6pmejHI04+ox8KVbIVO4ythI2L7NRvfhxW
M/oMqSq7K/lfWP50cCFjYIGPZXUfJjD/a4JxKbcCaa9XLkZiiPcZ8xxSCo6BE4PpW6JaC5qdbbXK
T3I5T3GKUkYbH9+K2fZJPiyV1Kc+/HBAtpApwnEFpSDcVc1rcyj7me0TJohe+Tz8epScF+nvxD4v
M4ts/iILtihduGhW8SflWuTNC75li3YcI/2grYYuROJpU85nHSs9RLbmUc/InmTcEAhVuEYnH2it
0CbX8DFVD9uWuOyN5jmC0hGLYkXwXRD07Gww8okaQ8Nj0N/krmzdhN5oQgkp3E128rKzfVfYy3JO
XYPSILqkhtDXeam5j9s50qAgp9nrNurzt7eFiVdphWigGSlT7yFWApw2Zu8a/4ECBfnfQL4ayXff
PussOVr+DfvTEMvZ2IsLkdwb+yM0w2lAlHr1cSiVf/pT7Gz/TDDCO+3d8HVniiAdAwirEuxjx8Pk
QanXsz2spxAP8Fle55VYQ6fFFWFglaT3Eok+PTVBD5UPeBtQ6gFcbZTHZtZUVXdjJyTSJlw2xzrb
gctl4/7IEyJcdf9IGfLFe5gCtRChU1gE9R3yOceIlYgZ2wy8TvClborrU8Iw9Gs28NjZKMmW2mas
/iWFjFhLnH21MJJ5kzajLgROn4Q5xigBjg9NOPGGk91rl2A7fSEftH5XHJWc1NLGiPZ1swyRd8AM
F5hJEhWcuT86q/5NHe2AlA2Lec41aDxzGmjnKKXr86HHlE6DUCTeFU84z5XQ/8czbHj1sxaPfWmt
+qb7P8wr2WYkAlAeAB56sEPNd/9sD1ElwiP568Xb93hAgr8KLfYERcCgf+38QMjHo5QbKHvpA7mr
923lh2MkA/umS/Lk7j2Man0QTF6ke2bBcNWs6x6eUnh73Dny7cyU0HdkZ5xWCgrvC0U8dq/IFQNv
ZacGekQqCvCdrErxoFv2Ay2z6S41sbVip+cIH3w1KoIOcFu5m07UnbkFo4Fis1HmUfAW6p7ZsYkV
CPWkOmZWVBrAd046bhTLvAdGrAM9jpvfa+f7iry07fsNMlev2bHFQ2b9/i9myCfrLvLY+UaSiFxc
EA3hC3Kc0+n5yw+XE/gK/YFTczfqylOX0CmjJcmrS+dB5pl5op3mZjSX6s+W70U0KxuwXBKGHx3j
C1EhOsTyI0s84h8m+Pg7nBRFP+qSZErpzOksW/46lMAFr4MS209ML65sG1m30IvLGXbytyD99Y9R
ZLIJVYlhvy045GbnZhtn8+XYU7a3xylauXrfUqUcN3Vh8orpwjQDSqbgWf3bDNCUYb6Deon1JAGr
haMe27/CklzV2ZNUocsSbC/yQnsHAzzrI1wjcs9U28p7llM9ndMo1zJAZ6F6YKUiITJJaaZ2Wv3u
nI9ImGgP4qunV7SU0fhODxRdR18TBscxMW+sHdswQ85VTpkS6EeBE1Hqqf1ih8cmGUvj2hNWCYf8
rK8pjGVu1Qy13/NW4dQobf1ouhvqX2ZQ5gYXqvcgTFifYW+r2iRLrOowZvHIMMiq+uMN6/cVBEva
Le1DpkHAGoPdqioHcwp8PCoY/TPxdHfIGQ/zXR0bDaK+DA/7XPJUIJ3koKLiZW5VUoXiTtowdy0J
Ng3kDStWhq3G/5JBtVsed+1Z6lNAGlv1BBco6RaO3G62bTkelZ1QHa1dSpts5oG19gvZexC7TYvx
n7n269dxsbrySKdcZ98dVWYTy+TihTbmYYuQOowbIBfOX7Fp/PjQSMuTJviXL3CI/ro051kKyPIq
RdfRj/H8cVU8ghdR5hN+DSrrLCLq6pB9vMOcKw/g+KCTDRxksIiFhlMr+7WLN7B+Uu0D5xXKTBX8
BRjMHm+vtYxfl/8VZ+WWA9z519esNtbpvbAogMfhhdUvUt5CWtWYigRLYjonz6ln+dzQI6jafz4+
sAwgXoj0zsALvXDjlx1XdRx1jLFhvh3sdGV+b3HLyGRHgK1Ne1LZq/QZ/phdFDBUQTvHtwdqVu/S
EqOJ/g84IUEbF5+prNVfQpvj1I5OoZhNBXK42s+gbAY1DhdqHclrGYiZzm8khyt7o7A46QZStXGb
dyhz0bnMTQALrJbYmJ33n9/zs5DSDJgBYwghEQdTtQ3oGgpKIQVMOFTtMJorgML/BSIAgUJInfTx
vznfHWBVIinzJZ2krBqiu/UOXVbOfxcHc5zA/SoFjDTY2wt1rNwkwspUnEc5WqM7pq9mwR8BWmRI
h1lF8kGtxdIlkv/zR5B1RlWQLUkclzZPzHmA3p3scHuJMZ47BM7/QPSNY6HduDgx380eKGiNsuGI
YZPot4L4tU5RAonec8WuAFTlfzF3363uwq1NYk+Hnjsf9+aIg59v/+yB6fzRtRgj2C0iXQpJJx2r
VP3eS5gHAWkPR7HMT2EHDcCMBGZgElmkoNMk8PLJYw7EuMiUlIKRVapT65Et22c7VTDGdV8E0hEM
hHYV9IbE0oCxvgRCyRVdk8MjQmbUyl1EZlmWAf6PmojOwh3Nfunhq9eT/lwUtn1KrWKH14f54vIm
dJAiXsWBIU2M1/RhELWu5Vsddq3F4/La5S79+QPJFC8erKlUVrEgm/pQ73oDkpaD0EqRsWrV0SJ8
pbNCKC6SK9TPxgmNTDpCAWB2OKhNSHvNAViMyAPVoHlQkkongqD9S83n2Xpxj+rUhTXiwav3CU57
5fdgRDmpOeP1Ewd2VuVsXpE8s4VjuczhspLZzUWq6nvfi5hoMa7BMZrCGJ+j56WkeJKceZ0bGoBP
rvfvMtdE1PihQQmtokMBIGfSop7GoWWcbQVmum7UuwtjF3qxylRt4VFIPLersRKibgwFrSPHhW0a
HtswRiT+iKLGEioMVI4NDUUpopZJJxUrjG2xvdnHt5BqyToVly7Sdhg5oKGQsgbHnAXdElFAuWPE
1hIE0X85UiuV1QmOVYAYkznG5Mgnw6RK/s9UUaZxb7zzns73JZhKr95p7XJRfY5l1RMxnhgsLXnW
d4AS8je9GQjsQPGVXW9nle8FVV4gMBE7/qu6HCMlZ9Psjm4GNMJbxsNok33IcRMcDL37bi+FtzxL
53PIBttzA4KS3qUcPPEPi+6fZz9RL16OhKOR8yLrh1d+rxaOWRmELzMXW+FRZITUwxfqKJ2X5OvK
3bwTqF3RMTAB+C9OEkdefD25KsBpfuvYgP8ELdoLCH52zMFh58Ivu/hlqOjW4lSyCPr9T9rbnSSo
o7PqxyMGzHJ7nIhKLkiyh7iNE9M1tDzEcL9VHQKXIDVgDFtj8Km5kQSy33gzBjJQfLtbsslRho6+
2wGaO3GElYaHmj0aOZq0S46VNPEDJLH3loYqZNfa1s5JGWrsc0YHia5A+3LY2spRBc1CktSF0Gzd
IbQWVm0zp1do6x8v9BG6U7KlgSu9UybPCnHT0gZI190Zsrfcvr/hrl8a6wujWizIrcpqOn2tnCcI
LWKRxpgcwXqCdkaBMItLvmq9WenE2y3WP9BkzlSWBarl5eKLcd+vBI9vQXq3ymoLYYgVqDGFtwfs
MOEjFnLCcibC2niMhHvbf2ixEO0DNxaLAFW+9U9HJ98jCHAweWuUiQ39lifHLMzvWvn6LgtBsvFX
xON53ZkoRmnggpgRZjRt1U4zIvEImuo0Sia3EFhyIyrUvWeeYAhxTLYAT5wEJQPQf8HJfZh6pvOF
+stDqW7D//Kf0hlRVycKZ3KZvxGEWQ8aw+75EjFwWWDL9djErW+2z7SsXeVF2ZGuAv0Zuti165Nh
oCOqka7gQGN1g77t6DmrFtyY72F9iK1bBqe/AFbnHWyq9MQ6ckKExOPyLs5lKbCzuVH9GQvQ618O
O1Gih54hp83D4aktDuOkNg5OIbN+Fd7q+hW26Lj0+xxWJufDuZV6nRVkHvES8ZPZZvAvEd2gIH5W
LFA1e2oaore172nfmzmbav2AMDsEmItrV0stbgAYnoMoZRy7HvvDjVzNmm0ZeOjv7vRQadreRQ8S
T5ruI1rsOxB5yZFE3UYySMiMYZ1uuptjLHva1fbOkQr+tki6gF4/O/bRYTMGU7DbVPBqHMMwvKJn
7akGHNwx4gsCfGZ4+7bH2yHniHrXffWHxtOQHQggl3zbGzy73AmqEKrYQN4IhAHsYxQ0vZ7ENXDL
Df+jd29ocJ8UqyaxBbuHZMKbjbN5YAJtDDFdF0k34SIAiPlGfgDPxW0YoVYX2GyfljC5QFKkEdYP
DayNIUYXqWvRVX15TwMgUDt+/IeTe6FetI5LYk5JKRpMXIbp5tKa0WKuLd2oFweSdrBEqVwvL3uZ
+V8IMv7rDbsivv5Oe+oZYecEoxOogXqM9Yw65/59gMoxAvQFVUjW03vcSscAHskwmu0AI+9POOhR
fCY+HxAacdhesVKTpKYvC2XKHx9Wn890uwI0S8WfXkVfq5onsBA6c5Z5dNV7dD/AHfC4BQydyQ0M
kYQe/b6VnoVO/g3MLMPr9XG7bqdDlpxXYQh86BiaXDJ1Lx8fZVneKTMXaGHAvyKDouge/JWKoIbX
8ActqSPZQKsKRqzw2IRlfMPw4A1H2t9JXAGAyHcEMqYLde+c0qpk/aTj1+UDOmyWJPowGHMPEG0h
Yya3aklFK3KqXayAIqdrh00FbnT/ocRxW6LpQ50YJO+Gpx/s5enNUN4pqMgpCHIqn9W+dgxwmPBc
wXb4pAJk6hD96X0y3VpgwVUa+SdJM2CaatkQid+m8Vm8m/PrmV1aJ3+E0SizwegOsyylWAfnWQlY
2aByVJZNSWqXUe1QdkXm7s3JIvgodWaZ3Zgx7C2f2/5hI20hm5gDWJAuUHK1gRQYWCF+WevB6hCs
MKhgi8/6H3GmYQZkfEJEir7RyNRLaBfHoYjd1I5Q6tTJ8wc7ieirinOaOwnYo38OKk8JhgM+hRXB
FG3zinFU6gFJuR3ze9qp5M12uof07DNgy4WWDsAYIK4VgDFmDGdAaoEXEQH4f4y9z1pKI5Jcwo0n
DjqvC3jlwMiTTBHogJEboczXZvi89Xz7j3aTiifPVwOCx2V9hKOJ+jsvz9F1BoPUnL7Rm1YDajPS
Jh3DgCBgmrdECQzyXlHnXgE3I5p15eBzMM/jJE1hpb1+BCtSg/O3zgTtRZlj62kQ0hjvnCZu8Kyp
JcI3bB+HwkGK3xCYY4k42k6pj9LDNQJhViZzyLQqZLSGX4RhjDTCaPwg/XJZ9fNVghJgFCWXf40/
JQz+Fg2pCOztD3fuEveIpKbQ+BC4Orn41NYSQKap/WIYd/8gTKXprR/qaQN5EvLPxwufimTPiD+v
sEKdLAEHtUVY23dGNDvww+4Nzz/MrSnjIixRs26e172tYqTWbwQGPgjvm5k0rJ7FCFpioSerRFNY
5NfDXD3mSdHMJBgPxFUzR2FJHpg8pLwgeP0oOKOTsigvJ9slY1uubprYvQwCKcLk3wY3bKelZeX6
WqBFUaG1BFn10loY/VNK9gaVWTL6qjSGoTmWnnm5KhV8ABSWJWaHXLQuaIz2oHgDYkBtdpAqj0y6
WsVy+sxhdAI1+uooYIPGQ0E1l6nM+rm7Iy1pQJoiCzpzZdpgxaceJVifRCmFweaJ7je2e49xsQzi
1RtcRRtTIYDZT+jCXAl3lpa0P5BzeWEkQRdOAU/wFzyXk4wP+D9c0o2AkUDBMh+zDLQm0zLAUOK0
oOf7QFcQKnvodG7oOMg/wRQy4tlghgUCRoa6gP25n5TqzVnovyj+O/zxcN5HS+gEC8oDQjYAj+IU
uS5bX50Bp6TeMqlo4kLWJIz7jgtqTgzIzYkImzN6wqw5zbqwnUgpBA9JGendaICwKl6xYevYuRYf
QWpcVR1rcbiTBdmDKKmUjjXeC7J7kJd18UkDElSJmgTNg7a/klJoxkWfJ4PDUpX1q0JoevKNgtDL
90HBF9/DQ7DRo6ka790td1Zv0MbHwt7DYFGjZvCyyktsoaukzu1yexu5rZj5taK2ymJww7ZSQozX
vja73yLAX6e7U5mLRtU0JELGs9VVyiT/Uh7HVHOmKIvgcyzRdToPELw+gSI+XB6KFxF/03VIsnRH
9Ej3lQU0/ZwsrlieAM0Meq6QEga9lZwZ4Grj1iyOZsNwtswTJkuQr5kQpZUgWKN5T+nzKuAyyQWN
PfuHn6TzedWqlA5Sy6JAeA2jdi337tdDH/TV2m7Zkiu1/gC1wEEEqkSoZOSLratp8ypisxLVfT1M
kgxiLZjhpdcNMOQHXcltQ95XqSC0LYqr6E41ZRgEIAoOosHIOsNeeaaSlnesGDzgltGKF8MJz8ti
iAIRmCcP8ZQMhC1lWiBv2rgCugI/ce++jtbyUantcH7P83G+bqg3pGyB2O7x+Z3v0nidDGf0e0r5
mp6ZjkRYA+UXpiFJA82AgaXkHuwr4GcDMN2u4yF/mPqDjMflnP6/+L+SHrHpIGUQLmGjJjyW40T+
IctaFvTbffuAD3lofduKM2cfeOl3qR+Zre57Jv5ZVu0XI3L3zJsbQfCojlN1L7hy8atJ6J4E+hlC
6EorIvg2RYlL7hzd2AT6AtoekF8yIEaX2/yC68APKJo1ibiI1JSBMcsGvII1DMtviDMweKZJd3JG
+cWHoT9tfzg1aivCiawh26dnIZfzaWL0YYFD8JwaTz6GRbQR1DupeIOVTISFbmBmOdLBoyAlK8ri
dWSrl3noAFNYdLKrG9vA42vJV9Js7eRRd6bqSLdfixtt6Jg0sUnf23zS0p68Kcy8E7L9CRjPhYto
IQEHxY5vyjuIb4rgMgKlfmlPxeu3uUG6OkGoPJ7YoC7G4c9UWndInRb5EVTIWzECdXD+PHXxNG58
pmQKToAWGcJP+NKcWyRumVqWqW+rLs7S1tQ+bPmXL5/p/Pwi0TAw+v4Q0XXQ/5NSux5/6jPbdHx+
szuf3OpeJ5lflBor6wD4h/dOotym61bWkPPhFnoQ1wbq9z811rgszTCZZTvjgKQA/uG7/zPqUTt7
hy9eHMHMpa384wNlAulH0JnkPiF6n2mMBftrQjBgUcY11yQ4sDKZGAI40TYSfCaI6EVYFRD5bFiU
j204tYi2Nh9Y1/ySq5KuJ63jXGBukTe/zP7N1bf9EDM6VeeE1RqHfsKjLFHLujFCgvwOvvVtXzgR
SXD2VD5Wm4AKh/TnoWApo8t8UQusDl6YxmYd0WF3zFDOl+Cw2jVpRiaIQQv/MknEsxDYlpfuwxTW
trdvV4qwAXhjoaPChnhbLh5Brn6y/iwdorZGHve3qcn2ktjcThB5j+ZDEXofLIxAWjm5sqn1rXsr
KCgPAJrFAjE9F2wP3VV42fRG+9X7Nbcvff2lBJ2x2CCCDis9IcSofdIIvpLN6AQ9Col2OU5ujV+f
e5vEapi7LEgpXwXJyVBFOg6nFA0ru4dibRZSVsdRWYwjMSB98oaGxEpPMu0Q2ux/XpbxhOG+/jrr
NYDVH82/X34sb/TcbnfloJAI2en1087VjpUexpB4Ld3IVNGNXPur6lUoYThWnrd5B3fb9RhW6HY9
foirkHRgSH0XIEVkdFTUrfNAKSV3RC/d/1Wm+xaUPWZhIxBUktTFywvfZcsc5tteJZfb8FQdeAZG
8RPvIL3OL/jHNlqTf6VwFBgkBK7V+q1oAPOPcR2PFNGbV08N+Ngs+N7vapA7W4jBeFKS23Y+M6w9
mgHs6It/6mrWh6563Uib2eJbAWre5iYf9899mroRbSFGfns+mUF6wX7EKBRDXJtp0WsIzat8NBuK
A4zbdhbHqhJuWsq71j/uCKKNN4CwUcFG5o3YOcYrxvJF45DAHOENirKCm6Rkw+rasUn3B8QvldA1
KZrp55tnFsL6StbwALofY4wCe4gC1FCCkAg6oE7NuMMc+ab4NV0T3kOmb/m/8f/+QBqrGno3vipH
R5unQPoxuyKSjKbJ1bWTI91tYyhAmTOTP2E7q2dSQ9OvioljswF7/3tIpwSkNzjIB7hlwPdZzTJj
RrAhFhyqNZxkQoxtNVVCrFOMVHZC1UkI72pO4GS2pM9amOxsxuYZe+fcqsH0yR+pzXZGnwPzMPCt
4U1gkCe1Zdkn5lMk4wbzBBDdsnS75XXWf4VgtsEUSz+SEo3kcRbMw0AhO3Y8wQaH+mYpO+ZvaQLs
EYwBbVUxCwNrBLnLx2Wqobq9BBT+nfm2sT3RXuL4gqX5TPKn/Dq8a1f59DEvp+6KMGxNZt1hKJ3P
X5mKPJDBiaSqiMknII5ZGn+tAV2PI78C/oDZbd670qTAINLW1zmk13NKWoB1nAfksOwkvQFIe3My
BbB9uaOo135OcwABBKAmvI5UDe4Xmmu4n2LXZHOCp5knT3AGbJSCe3mwOyg9GJ8a7SqPGN7HIggz
7t6hJXTrebpe6Hj1icxnF0ou62ab+znYxLZiqSBpgrGzg488AD8INhqR3xUa/FEPR91L2hMAK50i
bnV1uPNfuUMdFmVJVKR48aRue7Q9mtF7wOrE2gD8D/MA2343pAp4vK/Kf188Wp9+cJ6Th8UV2sca
oSPl6ANd5zrLk0A4Tyf0i7rBQ4DWoYiC6jUN8XqK04qyyay6h7VzWwoH1/LIzNS+6inj6ZwFDoVh
jEx2ys0+YUtV6l7APIuuSbOu1pDIdEjLccRuI7C5p+OHJmonXAdyZqWIc6bKkD6PUr+5SsS1268E
oFt8iinIxKrjA1fxlbZO5v++NJpQ+5+BEups4Q/ur6oRWTvIv/XEa30D+wKBsQQj1+d0BqS8+VnJ
9w21kiVApsVqgmt/lzfsXCyXpticYstg/mQ+POQcM0MRtsm8AOWENoy7kEGPA0LwtNdnXH+/FxpC
j/D71DH1vfKCXhLHaOENVSUgtl7DgcXWqoPPOBMn9yalAwA6pZm231BAChe/RdWpNN0QnC5JjOC4
IkH2H5xE+XZjaCBsEPuCOgN3990XvXoBsFt9nNoRcN+XK8KFrQBwR1fC7WxRMKgeCz95n4fe8WvM
BBy8HoAeAOeOzBRX7vMgER8gkaOnTSY51UwIqaiOAEN9xhi6u+3l/MFodAezw+OIRaWvvN1iUPhz
CToXDVA/igVWYaGEfpdR2PI/BY11q2fzSGyyGo946AHlFbsYbuuY37CpIJhQeNPrtyGDsg3iDXB7
7iAkqkiV1LLYcopGSc34hxC75oJs+WE7O0BgtzlqqIQtmVVEHeQA0PqnMi9h8xBoz+7sz+sbrKWP
d0z1ipOKSuG9HGip39Lgm+TCjE4s1JqpBUdd5fMJH7Imqsy691sWTkb7kzwOovLGl2kQujMvbUzW
ZGLfxFEAUhIO/dY+VVXHmCajANH9hp2vrJBqzkKhWAmrJUZW02FNRejJntnazmKBu5ZX+YhZpYBi
2DAozjKgOpXNOucn4JjG6re5b6qdcRlHJLJbThTFOOadLZYehCZ8QxMEnNPBQ33yuF8QduGLHcsa
0nqPcLqzjEJkTKMQ/2iUZwbr3Xk2TQ3S2DCNrigjLLmEoLBsEq57BKBBKQOYNBcIuVsZ7xdNWS4m
fVHFkjGEcy9vpNYBqQBYbDwCOpB0/Cy8i0mhG0YGso2V3Xkh3WXKCbl0AXZLrCWOLKsZ43oanio+
lrLoVqh9QeHfyOUl2HAJ+eWkfdn2Eg+0YjvkfQhqt8eE3RqUxmUXfTSDLvKDctrR/djN0ahwpouP
DzO3bhG4XMQr+wtiLOdPnn5gYovVqUeJ+YqUM90JeAP1XQbJrE3k3dpLxgCUGbXdwX+/zZLCuKtB
CMpq48LulZZYV3IjuG5afKChQAhiuDpbNuCCB5xAlu/SELxY5GuIOk6kfAnTg488SeQ97RJoBAmo
zbkoPfqHqHqM1aDAjLFZ48Tcx8LeJXguH/k8AZzbfmAD8B/R1867GaG+k9d5yVGUvEQKSoCgNDP5
skjSjMHj1rH4ol3Cd4IF2KUNqEY9iOSSb5aTf+soUsUK1xMwbxmobvoXQruUYLcfMChXNRWHBhyo
SyG4v1LnlNmhmr/aG/mBkKDEN7C2xxwXAsGcWnCMyms1U9xZx+HkpMXkuc459eu+/9sFnU91kBzL
Y5EztnOUPgbMDzt8im135y39B3cWf3u/bTSiH7JS8zZRu62CnXbkgxQN2dNUZIpRW2HAQWuAGxcJ
mt/p2iWJa+fuGFiYEsjDNqd5GnXnLp0dvlDzV11Epr2wTP6SopWCk9LcCIHmxyRGG92BTlkt2VLc
GRAtXODTInScTHgwbwv5PIV9rqxI8N43ZO1/6qgoddsaXye/4aO2zdC9a3eIsl8NxFX8atc1QrIH
PFb6RpfpcGaJe0wcL/e/5TUzmPLIZ9nlaJBVW3dRxLW0hwEp+AGPcvggyXS5ambnU1HB2GAJ1RmZ
2thw4951A57fNGZr2bXYddS+uxhbwJIcjuO1F/Ko9PjRsfwtkqyC/UoYFb0h5DQ+E1NtqEp9Yp8K
mh9EYN8pWbxm/+eh44Uru7+7ZQ65Iwps3RlI0HaL6OFBGtPshBmkUwZapRBemwXhiC3RWPtIZ4Nx
eqydiHVtyDKPzk9d2DTUMBTijkIFIMDWGoQXS7+2c4ShAa2uAaNeWoQDWnSpCDiq0RXuyUwYJTOM
9gyJxzLuuO0tyU5RiCsCQjhbU3gyqCqcdN9QWJlEDSZWbdG8SBLNr+oBgcr35TH9SA0QvSJLBxG8
96Pd2JQMQYqSpEYLm534yMi5E7MLDjrlUSZLuUrHw3W7+Gx5feXBxB2tUiUCx/8rOruyC95ANw+Q
whRfB3hFEgYJ41LmukFt4BroqNr6ehMVd4qum6c8Tho4QNT7ijD89lCbqFhrlKutbSNn3YDqR2Rl
rIEGtZp4eDUVS1kS/49tSSawttx/2uTvRWvYnzSIs/Dqr1OruzNW5PoHvMM7nS68TWgoMDiuyw89
WoQ0ZxIGZfsgLvOUyjxUOIvP0xOTnlbfBLfso4EzT2KsAuEE5Dsn10Yk6VIu2JALo6DbTDopNCLZ
fgasPOwSNDkLARJxT44z1nXeWlR3zjmMOfmiThxH3nL5rx+Oor2ZfFkFSrfLMdrjoBXD1mZQsMMh
It9Oy1qVMoYd6eG4wD9C2hvLLWmS2fjUnRij9Wsjo7B3bv7HcCkhxPD68+sM+iVsRz8f1SoT/En9
joV9lUh76MyU/1nmZEDQ2coquuqmqhNLhQuoIDK9IfcjI2z+bT7w3XeidK1DUuOdfVVGOH/h0+OL
nedGVf8mXK6/25XA5X7IxNbBqgOEkeNTjdo8KhJYmMMUVrR3ncuf5oeWL3EpWMDfxlbkSb4jxmsI
6fENMpJ1EfosMquKMy2bo5U8nVkyBTtOgkE3lnOkMaOksxshPqHV4WxxTAEofSsA4nPLnfkqNI6q
14M7bLbHUzsiW0d9oRrMsbIi0X0UnkJ2PNl9CxtRgt3QMkfZQi2V8zGwRwocypu/SUOd74hlZGCU
dvA/X1GIjJmZBodndPtH+oHjud4dAgWOF62EX89fROEEe4Igz9UF9MaEbtg9AH7h3rEajIoSmrcq
mwlvGbaNVFSvl141pfjjxmMCyvZGoOMim3i2iZu23Znad0EWrEK5HXQHJhfon/vUoBIORkDT+i0r
CFw9CJWC4T6CFNoDfkJ+ZzBdwoCC6sKoa5L3IC4yrGn5vpN/HUYaLWyB9MjFquv9u2VKpWCrtdme
F8Jg9HMYlk064lTLqmZ0WmXvf8bKS1YcakAHB1RmJWU1uF0kzoF2zTinJeueWNIJ39lEYFamkBjO
B0xGRAZLBm9kiPNEgQIebFWlNwDmcDfjJfzBrZjjV4JgpGxewk0PqYZhl0GHpHygCoGOnYEyCg1h
N9DK1wvo29hrJdHsF9CsdZUovlNjSb1xWwZ76mUVdN0YVKnwAiIGoL5zGcHGwdk2EiE5iGKRoEWF
GsqmRHarGsTKwgHFVXTdlCzG9roQmAkzmpemK6tAeExfwV75PvwSRAnHILJOG4kVmMu0mR+Zuv+m
LnDaqW6GTE0mL6mMKDdbJVPP91+7uJ+sKiJ9iR1jO2wAXjOYZOIGAGnrB626SzLpRULud6tZL4Mx
67W95diXEXllVqAL/EthNe1IIWg0mRU96YflsSjgJJ1gtSQddTaBQRzvEpGr/PLBiWxs7rmQ20ZN
hJqH2RLf9j0GhmRYMg/rdUc21Uq29fwIcW0Cl4V3I9CBcNy0jj+rxcIS5JLQK2I4L90tYGxN59Mr
OPgTYd82m4COUWP0yR9NFCKR4sgbadQ7a8UHWxiujNKAIw2AUKUAGikrxyFE/NDMxIcyvQycXoVU
3s6Hz83GBVddziJwDRD+EltkxO1vO1LR2DMT+Qi+pypzVoRHETNAFEM+yYmcRg7VH683ZlD2FJDG
jTDB/wEzwH/1uMngL5cpZSY2nJdA35achtD7BuvUcBO02YZCy5j0OZPI1AHlSnQ0pmFHPYUyxo2y
iIwI0BVMZXu9jBI+iY/qW7JFNEavqt8rXNOdPzWsIayQHcWCcBEW26sDCGz2ZjkYPL96st3yEaBs
FW0NAhWhAclIhh9+1MVa7wCFCw6Co7kWKlV4CY5bB2PNVOfIKKgq65bRUBDymqjlcSRKdTOQbdzt
J0Flw3NL0s2sBWfM/iOu8nXPAMuI//weApCDQMgdLfwDqLQrF3yTjDFc5Kf7a6WgWltCbBe5a0xH
aiciQA9st/0SI12w7q7kMcDQOVkn4AIqyrguZKFTClfLcKug1BUuVEPKBqaJc0FFy3eU92zLKoPC
uahuUmRG+YFlUtzJ1RndVbAiINVW1E+79pu7KQE4As3Icc8sckm96ujjm9LPTM0ifXOEHhWkb1LD
TrTZ+syCyTXpKa9iicKaL3q2PM91E95lmzrJCXEqJIt+DcusFWHvrcqYhhaMdNORN+eoOtYvPQ5i
4pQLRgia3cyVLgrMNs2CyGuvcATeMoD+FkhJG7j23fsmkvTZQjFzmfWdmpq3OZRA9RSoqp6x8tzl
SF9rSXmvRRKUHE8h5WIJ23P0aXV5jlSHuxSmjt1TbN35zrYrXz2heIRvuUxuCuTb1RPbDgF8sQhL
bOl3iseT4WWDFU6WTxbed/fPBNqIra/RSuXh+HL+Pa1IR61ghQoQ3qivvkCDvBoqiXPEx9QHba1m
3ty3tJt21pmOaBx5Bh20oiaLX9UW8dQ182VOolV5qySdINrB78PLCLrmFYyAYdEZToNHQC34SZoQ
VFnxxF6mMR6Rkp/HWDHbmydGEx4iNdNMnwwOhz8ODmpCpELo7Ms0TWBGarwcGse5Zfx8Rcs3xL1Y
PXcXaFV7I8COIo94Yw7Wu/k+OwswdNdPzObeOhymoo+4BsWQWNRUjo+ptX8dLnURQQbS1ZWIfS7R
xKHqt58DRlpYqxMSHK20ofLiFS3prPBXud+ej7mEibC0CsB8Who7YcaxD9xyE5KNCKzNgGhS6iGI
rfZCRK4bpwuRD7GSVQ/Z2fiJmMVHv74av3DqsO10U1Hy8Q1NdZYA2iNrvIp1WKdIccMp8oBSPs19
iXzAj6pHqNqk2g68h+vFqrQBneWZ2eQfnAV+TK8i/XAEfl8TJLuUMqwgsaFnfoqelK9LPNT1ujcO
+RVuO+EH6cqJy4gNMw9WaGc5/2ysssSNegTK+qETcA5RCgiXbr16YURtPaTYtoNx8OJhOi20XJpU
izuyRmdY7gd3RhM/nRvfTV+4NAw9h7j+y8CJYGYVz5Ho20yqvw+2OojHHR6z0BdVfbhTH1YzVSTs
c8ToixOA5pIPjsm7LhQOljAN+0pzPpnSH/fDKR/vq+LrWicnLEMJQaXdXv1fM/McYV+gtL71hNkj
IwWekSrRTGuHBAx1ecByiNYcBGN6/DxjmroCONzUISloruQhd+r2k2WW96vps+4HjJuOecvNuXOe
5JgwYueJ/PRhXb7Rzx6hjON9vPwdXpsGiQr9ix+Dr5L+pJzcLvbJpaF6m6jxO23dBHuJx3Qh0nCj
rDCdu2h4Omzqk86w57ckIISVtcCLsvpbwgYJq/G0HEnOOz9gS83Igp5OIdmRV9trL2NGxyMKLjVF
RXkvWAeIJZmE7q+LZBSp8C/ivMUh2O4uGEzxKUU7kgFiQSxPTiz3mLFrGX3xzX8qFSn7e51EtuXU
mVYAeSqi5eGnyzkxmp8gk1zu4FAn57HRoIHnTPD/gFzFglh9HFDzSL3FlRFEoX0GLpbV8T0Eq31t
HkFhJW+xD8bmxt4B4rlkGh5Gc20EyKc099+4UXn0O0W3DgSxpsTFfoZ9A7xOYPfNtMvprXIwDK8O
r3A3qHK7Xj9o/B7r7C/6DJWTyZO8SU5CPkdrArfYR6RLO3p+B2xyV6vG2eRafu8hI7A552F8mc7W
4JkjpFn5oCylSq8fFFVgo7beJcqS6ljt8tKfK0mmKfqcYNOkS6piBrf3/2EpkNByGEYD5meUxBEw
LN7viNP0dRg6G1YHRtKbsLto9ivhNkxbxy+FXC9fVaP7Rb9vvAf7Rq79GPkWqzNcNBKTuTAj6hN6
TiVC11IpJ8Z40hN9hxpx0X0kCio2Bodwn57GAMn2p45hZmR0xcjtv9plNkLQ60nSYOGecT96QSbo
04UaFUWGbt7WMfvfwKc5SaElUlKqIRdOLhZgq4aYRU3jejy9Lu0D9olGqPN63qLcPHviBQgJTK3Z
1qB4nQ0rD3R26DXU7PLxE81Bg912aYlpxsa15Xa8d9XGmN3TbVyr+XJBepBOQFM87DL2UcXNihtf
Xwr6H//EdwbDtaxidGhYBPnnAMdG8Jxs0wvKoLE4kivzSs4YxCEgVvVs+8kC/E1FUJlfdhG1vHm9
ELlLyUVM8DXAUTS3SZv2lzauTrF7QzR9Yd1Fj3e/tH+GsgvgtN9+qr4Qzmifu26ov/VpgRPY6ApO
GNNejRlAiswVJNKwgtoIJKHgVHXdMn/7nvYW6VWjvT+T7SVmGJPLlWL7fH1LhSFPVdgFcWyftTA5
9uLwt65MJqDDKSxp20huOw6/eyJXNJG5QIAP27THGq2IgDrqegMxCzmHQZsAL236cooLKaa3QtSC
rJQ/gJ2dBhOEq42H+zAMZoFdlfSeOrV1zdBDDN4ar6RSyj5gdkxYTHjVS+iFn0luUp1hx4sixhfu
kefQ6jtEM7sRG3DFFQxjM8neIw/F1RyKCzow8OwVCfC6xpELM9sMjLmcFG3DIu6XJ0nOqNSnl9/t
+IbR7rehNyc5n+E4OmKqK3NOAQWUeXGCLJzswv40Wa/E14cTk1b5xA0ydA0QPLfH0mNifz9bzfGm
47jIa4i5CMuHzjkcLz+10CZN3UDQbIOPHFZHw7wZdwCfZV6WX4yujNM07OXFccx+nLCjRwJWeZJU
TEglkkJTwpIK6uRVlwfIkYMWsLeoYS7w24xEkolgsyG+BeGAPyn8l9yqd6oyofeowBqWHSMxdwrq
WY9JKs3uyA2sypGxVzfu3GLEiN8f6c2H2aIPen6ei7MWcu1Tg+0p8Zv/dwr/Og3vc9XoCRss1tDf
nPqqMabhm5P6qMabs/HxltK9jsh1IcjFRU6kJD7Y35eNAPEnCfJTd04evpOdN0mpjP3dHklle6Yr
phEasT98wP99a4uv8XWZESxUbI+vUUbj/X/YNy/dwcVgPKOTjS3pb/gPPUr3f88Y4Bk/0bqsUl+n
syf9tc2lMMfEzswFkC/iLBTZ0tjGlLBHKJ2ctQ6b/9bMJKeMSIi4PrpoyBd9raJ3xowP+D89k4wk
F4a5hVLzE3dcKmqWQ6m2yUqHej+mr8uyX2dqU/gYtTxr367b6BRZ0e0tKacLAdQuSBou8L0Qio3c
goFkyX/qlQr+JxIEA3Qqkq7eDuw2IxW08qfL73apRcarS5WyVtWw8v7I1PlxUGzwoGHt3h4Oe+xq
ZZHs6CaYlZe8xhmRd24j/dCg1orEnOyLpy7zw3h6gkTo+E+6eBeGSWzuK9s5JQxN9bH1gLpJGUe7
4lNwEVI8vrvemdXbyMVGzbr7oC0QppI04kQRMsVaBSAoXo20f14UqBACe+0NGi8nyzTukg2+WFsB
fte7MHenDOJENDpq2/JKqVQlCXwhF57vM7URxbnDwX3t6mGw5YS/3MFSFtVFfHmWlcn4uWjCfxvT
tsca3IzX3CHMC18bgz0lIFkwbPWOiIxobDed7OdIbyOFtVVTgN+Q2jpWcqx/UlIsTrf/pnMHnb5j
r80aJxbcnIZl/DfI3sqrxpPr4Fz4D8/QUSHc4pKASA4FT0I0yP3+CSsqcNZxmdegSCrI5CeztjPr
iwXrlDmSDE7yOHwXqmRJ6s/iBHJkPg+I+1NuXYTx+LvV+edIAElib0cPdGF75zeu8UepX+v332LQ
quPKgZWuyScXUrG4xPmKLGuw0h55VyYq7bmUFkQZwtLvIb9FVnujgLe8E9ulQKbMaDsH4cuJWgCJ
gjZMVk+3YV1aLftr5tOobO9PPpYOCiZvvhyFyREVhSg6AS4Es3nMh/XXG1tbgYJJouTSMrIlxt4h
VXeOyaMdtlst3bckKkqctOQTc9epCh6/01dI0Vu5NLCys854lZYYKN4M1x9WuChxCGplSAIx6Jp5
E6O1IcmUdCxt85jUTQzPh0h3ZVdiacJPMo/XhfBAEzvvRsquleG2BgpJ9/HyzqWThb/jLWDOwCRS
L9sIgBG5EPP3w/vVPeORmxnc7H6lohbY13T2RO7WiUT+hDM7OXSls036y8XVGBNefKx4gIKqc1Mw
qNzNiOKmeMGN/UCVmh1rSojwIRXoPOZpgngYj+l/Je1AsJEsVc06VS6QrFHLnaIsb2ODRZlzqaj6
STdx588TissIJTYh9LU1Rjq5pA1BUPtBK9MBjnvt6vHXbMqVQ/WZi6kIdHpToCKVUntkJ6EoZAXa
UiIKR6nd92di7Gi70LjJNVCMPt/ovmS8focD6OfpNW4wTUOCncjB/3EZWYbFn6BKu9A7/Jx4LTEN
OfL0pSFfIBGh5llMuWHN+6q26eFZkCU4w0x9Q9qaz3EQOzn+Iq2JHrx0Ppgz2Gs26L1bYUZe6zL7
QxP8tsiohb3MgHSfY+ghns70qvODHG7FjKmuISmO06xHFksUO5JZUHndnC1u3194t6CttGhn9zVX
qYiEQ5Z3X/LtEzoQQR3PnRmSfUcuzU9u/fuhPJJh9/JijW+sGOAFQoZ6yvioWnTLzZa67JMBtfGg
XrBLaGuuoVsu/raADS52G+Iyqqp9ONfo0XW32r3n6eMdEBMxABHUjU+jg0DjZ/wscxciKBLnsB5E
BeEvVnUoLbkhaKk6LhJjPd5TcAPTIlcdetkFTdCr9trYUrBYgKW+1+1dHgKvidCSHEynyV7qFnT6
B308zakgZDWZ4NYgiswrQ3X4owhh/6+rpNPT2cNmgvj++CSlp6JFPpyuwueTp6Toh9hS1zxS5RV3
PgPjH27q0AbVGze6MoFm6rcFdsDhC81eF5uY72cZirNklHQjresHov0MKeQyW38lstQZ8kB2mpn+
EWeSDst4bJRrrnhWjNjY8rJMks6ZQoOJF8xNeeU+x7OGih2LyJDTatcQEOhNalkYocRGpb35oJoi
+rj4mMCvw04fjYrdbwXyW4UCbZ1UnxpeNWLCZ7z1YEg9B5IY+NxuVRd8HWD941q/pMVQtnSesvpL
TZE9WKtdUCfvCvpsaWwlFe1eqnhx4r/8+zbGOgHlXpBwEAq2X3nIpf24WWNQWjvgGWKqpIh00YFz
KVUNQGsXT01VmBeSq3Q683Q0iAD9PpMex+DsjmHVhQtmkO+U/nHSDt3/GC1ueL05MlO8ludY/cXC
pFR7zF+rCpNYpwV3AdVjo1QLUJid8CtjTi8Uw5ImaGWKWgVOpOIQyP7W0zR460vJUrasYs0M2LoY
uxmhPRKBV3ABqutnFqJOUQfdnNqCIhzYEX6PmV1sPTyrnppZrwjvqwBOyy/ePXF6q/IkOvB6iUHG
wj25nvvQjJnYucqEd760RjcSAhO9kEDIQ9umsZQCECnglp1tzh99mq2wFZqxW7iFtOTITTzsvq9t
f9vMbR9YlN6y1r/PCsfvVopbdRYL/mct3wD572adbrUnikdHGrOojAGpvs0TNBTXGBFbiHHFO53y
amFptbck9uRukOCLgMb4vqNoKnf4MY0g1/wlI8HxDCmKYdTEKRye9IbjyYf5uPPyLCzolTOsk+zC
emgpgaTrNsoTTfv6EH/DXv4wnXlGq4ffGJQsOcNgRh7KwA4zSqSvKUYVnD24CF/gl/O9s5si8T2I
PH7UIoBWAGZ2rcHbAVrLLO0HL3qnEJtTBIYcgmzjq/8K0J3QlIUJ61n0GtlHGCfD0l2tKqONnWRi
BteEavuH72BkKj2zdVNxQiyU3W0Ou+4SzpJdS3MVdcwxjAat+mNkiHHp9uqpsvTVU2AVgR4Ip9VH
1YTqWEWBl2F3PKXJrjq5Ev8mLvz6Sizaku6wNNHENiz10ggQory169fW5x9gXWwRl/yrsK8M6BNz
exLbJG4zom4I8JtIlLa3G7zOaFxqH05vHvmpebTspUezDqztc1yy6hL7jB+8cx0i/SQ8rNWlCdK1
nLNdoFoMTsgh46GeoSrTBxHxyfdUgYpW9gVh0fh8we2pv0HeKcKlvSgVZ47HddZb8aN/njQq9R0r
Vu77TKfPCLXiLR3l94J7AZF4f8JCKnSzmXYQMFA26EAGcWeNg4p20EipQGpQXwG4NoVLjDe8nJ1+
S53ycmp4/7baZ3Vuo1TwrkpnxUfA0J02H6oODbq0DcUOPHcahJtWmJlnxzLBJBm6TIANU9AJs4nR
0YoINX3PyoocXPcKIJjvW2fCR4tu0BYqu0ggwhjC3A/4AHcDr5cw17KPc852KpNg9zkSNbANV6CR
vGz8/kfJjkBwuP2Ukr6HPfpmPwGDT3bF6pTvO38Gdj/JWTuPkNq9rjt7MgQbSdB67TYMFiW5MgpH
TxvIbftMN+CGwWqzio06f3psrXGgkkn+ppZ/O7r6QJ5skvLCYdKCny7qDqBObxqpgeUqZjO/QJ32
sovyfp9/HlW4HB3CM55VOc0a/tTe5XYo487/D0W+siVTSiwLP5B31gU0yK7yP8PfKrfuiy80HLoZ
a/k0U0F4ZdQdx2DrD8wb+2iLL8mHG3OrKC5BSfnT69cC54rUqXG4oF0FHPEDMSGGssJhZ+YEgX3b
lgObgH4A7B7XlpOgZiXmPu7mbqneCuiaRzq6dfb7rHWyjGbeGWE0oJCvQ1YAwKyevDXas+dFXRiy
nfqAyHiiDW4dsKjFTPV2pTuHcAoIfh88QJvy1UJv70OAZXta/Ji6OjoizLF0A7XsedPoepF+HIwX
+f64CKlLKrV/rcQ8y83amlpAQ5GVmnQC7GLoAEqiC26JHEa6FMdus/sJqikA6XXiGHEs9sX2cX6R
BtM6G4c5F6h/bP9RVcgJvTfthpjif00S8LjCsMS2FncP3SpFnR1GMkrwZx8ASz92qOmJUzajqNzL
4g3SeikqqVX5Q426eIIfQPIUNc8iAUz4GANxw7u7z8svqNBckWm4E6caYrjIsNtj0T8KccnHDe+5
GY2SiwZHppmRfxg2fCVTPhnLJ6WR5op3YpH96XhVagTyClEF0huuNfY+2O0R1wkrm3oBRY/oqGxy
80FC0gFczyWEockyXLZWnt6NKNBtdD/sGv2GhX/f7EVNTQ21/11RvF/kdBILRLGNH2mRhLh1DcLX
wIPBts25nMAZor4habQ7RWBx5phuIzGqTGWVLMWB1wzG8f6Q+PGteqmr8+yx08WPI+tA2sWTrhZl
eeastzXRWefyM/hd/rEwGfckEneoXNezD8iZjPfBOmcF4Y7nnntf7CQXWbwJvaGVoBEIUUznAj5r
RUVXfLET7PprzwiS1+SmE4VASCNKtCddSgWAjwHSSPxUOmJJti64GJyZAM5pPH2o7wsr7Cg/1/Tp
qtFbMObC3JgujT6qjfhYU3N5XDgtn89vwpzLU6vg+EKuO0E+IKF2nznvrHt3DsPUI+8vhAMKQhsc
DWcZ95XXZd6bYE1MW26OCU0UqATB7YkOfy2IzQi1GJUzRUdO6ZgO72TnvJnh90J84+45YH2vIZWv
Kcm4DTcH4eFXcjShJqTMtunsHVvsxcmamTpTjt+jFeHWhmbxXyKDVPqDnILAWQvbzJtKq0Uy8O8G
yS/pv+LrdMthyJvupYfaK4Aet0bq/R1KFGTJbc4oRhouATNIpnUJWGjVt6mZ100bPzuKTjwPJPm6
t8FiGqu8PEtmerJ9gu3qFoV23lvELpRcQlgyqvymrf7izbmY/165aWDfggCJgUYUlUEWQzqz49Ew
RQ+YIcJZLXFIt3ZC4cZAVJToQvKSjtfai2iAgO8M/pKzcMqhcHJL8oYM00DX72m6NrCyidwB9LfH
vNDkPH95/kku5LdE2Liirpd8JnFVfepdA2LeCXYdIdCnJ54ETLxO6hw8Mdr4kaku0GFnk0/25egp
UZgcb7BG4bCeBqW19iNY79XIDzEnoMi5k8Bw0QBTpdKiXiJDmZ8Jn4PimsU+GlcbIMNoMBLZC1Sy
tq4pGQacTgVRLxfWPc5yPsXSM+Cl5zuy6vF7Lou3Myu7n91+oninHupCp5poGHQmhjbLhx23rw5Z
Nj2gQqQiMxIgJ/UTt1AMhWuYu4KyXOezg8CFRWXOwX+4bbTAWQQ6vvxLwy6dvBlobiNjN1PEcSNX
dTipcrHeX/jy9Y50JqNkU6Q69O3Z1YLDzq4adB5cieghSKdcCrRa7xv+du5f+YJpM8kXRqIUDB19
c1zfrYe/kRoEBLaV5uUvUbI1oz0q5bXd4gfTIwAMonPGlgF0L/QLT8RUylHDbIP0qKndGI1fSVPd
H4PLj9od/SDim4/VJydU2h7OxYcky7AI6xZzXl4UogRebLQ0y3v5joLgKTYXpEbfdrHlr+j4jpSe
IzakIf7W/ffm8bmBHDZu/vqREFFAkQg5Y2DeEWjn3Z6UuUXiN2wnyA1qICm/OpDFlOvEiuHAOeQ4
hc3ZvuWpvYjy96mBJ/kDKOt4IWJOM+wGngqVJZTpQvfyaQVaqnuwctquiFkJD2ciDVyk5QNv02Fs
+f/8WLXGCgFVK5lvCP68JddFybJcWtblEC7Np7UegrtNBoG4jgnx8Y1ALLfrkBYaM/0LRFNjXVeX
VfZHV5LKMLjCFNvay0emh3aci28saNPXpLF8U0BPknWKhAUkMhBxmRFw/quW/1eHDWLoeN0ZLem8
31d5TzX8ABBktJu9nbSUCo6ZYl3+/5dnkIeOAYcD1UHOUfoklB3VOvAXWyVuscsVVQzbPmuwHwDM
/x4x6rv0cD9UdAEBL7fO8gPbFzAkLplldzWAjDjlyLS+2fVWNCLA4zD5q99lZehBtl8YxI5orCns
W2er7UtVL4gXTNJXd3FRq94G3mYotWqPLLjLvK3kD4JuYvk2TzCibqb1ZpVg2S9d9UagdPGnEfWB
HkmHXITw8Vro9Rz+bv45bXy/RaDfD3RwEtm0r6eSfETyDiXPXlRnehJdKJFTrPBNTBlhs5bSguNT
+EzLwI7FcCO8KeGDwkP3hwVr2Ct6nEU4Gqqes+omX2yfFMvBwM1Y7e9KsqdSR6F15fLBctuokDCp
fN0Mf4WWZxSoCrJyoUAmZikGnCxxKBVn2YRQ6ywxzA3qidHnEGfq3ak+lBfZG1YQZWf6GHovGF8J
pVn6DoCz0NZ9+V3pD7eRUtE7iZVuMgqRDHM36Zu2XmKlro1DvYzMM9v3l/R+7ULp0/aqo0vKcuB2
bEU7DR4pSLoKNOzeMMmFWdwYEtK3/j6TlevTig9BST6RJ9SCAQSBTsVfd72J2QdGm4mmC8ocE7ME
8RAYIgMqCAVUr7mYtcAEs3tU1Am7xLURhFEhI57Izue9UxBsFEfku7fCr6jD5NaEurNUkGbPeWp3
FNBd9xdjD75Bf3uNRMQZzu/tp1UskRWqmd1ymtAH/zDBTu/m7fnwJSFHxmju2IZsFp+cJAHuKTGp
ciBMI+SQDWJRq6vrR0BdsW6OSTEmx+t24MJ9qeUv/YBZdqPobHbTIgSeot6yIetybzRYInU42SLK
kHQ4Si7aRKxmf68LEhlXluEnDMa4W/FA6ADsJ3m4Rk1aaSfDuScxxweKYRVHODVei23Upf7aqfeQ
7QBjV6EGHaOsJ+KQfi4DO2ojMcqMwHTbCy+cEreMBc3doypfyx0kHEyG8RNQfPTE4xQ/E3kHLlDn
vE8ZFWlxX/pRXlfChzIGoqChvFf8IIVV2XbBIFOArl7HZ5rlVg5pa733MRtBM/l/zCmPSm90LxI8
lDjd1aDB2mTNy/2gJEXeac2dPWUrfvu6Hvih8gKk9IyQ/n7WoRc8RKwrU3gmPr2KDWs2/MQsKo5F
joMV+8otRNJ5Ci4qjOsxQpjbypZarieD/7hBLQjGEWdwQOQmCf4HDv83G83Pt25hnJ5q3n8xWy8G
wTCSCmziKYx1sMxgqP/w9UHZmIElXSLo7mfH98t35+hXeQD+fRZP43wAVcxiwl0/2p2X3+Ez72+h
UB20Px/S5q/jR/mamulZdlm1MLRSHpyQ4IfnHDUczuAOnxfEFfom9PzCb6OzB26UDtJfJlHsngbB
LEBH4YfHLUjPgpzFB/p+Ia3ceb0BVBoIx+xySdpegMYwEZWQreRRjAOAXoxnEzwtnEdhEE4h0G19
bs8iGb18Qv8qGs6M6gpGtqZXxsePPc2+qZV7OqSEGEEiIp+Qr01PmWI0RjytRyx+96ABo9OTnBJe
bU3e2aLtxzgzcHwSnDyNDw+HefsKz5SZdvVMu1E5/ite4wiyz0ib/GxQOF94HTDKehVlGYdpHb9J
4SJ0RRcLNCLQapKZpNQxglJVKdEoFeIAcngTvXza5zWY+P1kPCBk0/yh64vByhRvZNQEm3rZ2FG+
6DE6tYQMUBHaLMsyxBCRLHRL38ZwpI7pAKdyQU+fDoqnsrd5ITGzO1bnekCf3mOSygpZZZVHzScn
wuVps5Bl+uEiZ+i5LOvNisFZdBYOKPMKKQCLD5+gSV0gfB+IUhgbx8YXibXpUm/kRykWfTD2Pd1K
KWr0swHMnyjbidd2dUZ4+7ab/ows/SLslWvW4fL99IzDj21yUCOw7ypbP61VkN6zSmxzDp0O3gtp
2efKbVBQJwI+NAawWGFinzfyB1Z9BrGTVs6C5HtKKOOJ+fzNCKvXUD0hBZzdoG8IJ9U/V1825teW
brfOzUjHE38si7NH48JjqdICshm5kg+CeZ2Nnfe8sv6+tPSzyasjRPFsIPWDNX4bYnAYQQL1YJ22
PSMl7NvUeKJRI4wmrGq6i2b2jQtwxdBOu2ik/Md1hPzr7WoPEHqD6QzGHdUJ95dlalG31wjXdEgp
UBgslDYLZChD7nuxn9BIhNFa+NJKD9b3WxuCBAp/lz9tZhgPLceFfgsGCutBEFYYaZ+Y7mFQ4I0e
zMLxofmx0tvFdk+EaEmD3rgFTJ8l4RtgSGQx1igwPAOyLW5FesT5hH/YcAJ8kAG9ibh0bxU0yD6c
MqEz3WsWRUkotjnQsC+79SrRFbzOHxL/8jLZCj3OUBH4UMh06SIZh7aze3JFdC2VaPuTqHDIzw21
A2tUJENj+w99VNnTsW2RcVBZ2WWDRh346Nch9WBrWu+xJ9Dzwr5ZJn8I2Y2zzZmdgDsRbJokple4
Bc0MlwUmRcjzkUtAthSP80mEOCdyJXFCkDQt5WAVME3FwRPAKdaMh05HURx+AqsQHtxYaUzeYXwy
Wo/ufRR/PDh6zJt5TYz9MJIPzDcoLWwBkjo6nezizH7TlQyQ3P8laRxkgDD6BPcuBmW3/syZS2v6
FH4Osn3GfCASR88BpdIQ+6JbeM8MEkB21T95K6cRkVnwlWO9Y4o4NziyQ/KSxTyG7rFk9NaIK3S0
WFwpOg76tsUqH+E8h9UAWnpzGY+D4DuPHSNax2nQzL/FLekM4nl6knw5rXhF0VdXtG3PmVO2Z7r9
c86ahVZZFPcpt8wAfsA+ibdZlYxJexBzkUWJo88loVMgKkJFty7e0U/PMv1M0sH3f3gTumBpNuZP
9c6oqOVonTgVuJGEu6no1XH3Ax4Inye2ougEBTtxUqwliVtCU6nTOyFeXoaeg/T0XjP0bRquJNb2
RPv6jDEElJ4tfzKX8oh2fGvx6smMb+3xWoM6vzKVDwWdY//BNhFSDcMuQ46qPh0jcUhx8KNYlENa
CzzQOT12LMVuzd6qzHqAAhK2vSHhnQuyaWY9tJ1eky9SGU8x8BIivm/ikCSq6QUtm+nmctMtm1Kg
BTVF3zRnsGYqPZr1GhTXC6kjP9VyS/OA4tm1VCE8lHGd0G80piMJrNVMr6uciI3Gw3pZgfraAwmc
DbHPqWLkcy+fxT0lRX/NhRU0IahI94fNcx/OSw3wUI5KqE1dtJC+4Z4z7mEvVFDooEt7XRlj5n1V
za7gXXqLTysORaWk4eSgJvonz8q9LrAw23ZnPV4GVtbsCSZfG3AsoLUACb92BuMaq1WeauM8rOvo
o3Sl/WB13BFyhIPLLBfi/GZsVp4SEMVAykPkZ3jDSEDOdHeQrXFU6sPmNwfh9JKUf4r8cR2ADW71
6Uv9YmANjuecA45grjMWLVzXTvWfL923G4XoFWUgeA5kUtYP6n/rTlOwEzpyaO3XwWDJtVJ3EWyk
JUtf+aRspiCRdM76xkdynhCariIKyRpkEFLsxrgHMi0QFr44QRA76VnOsW+QctkHtDP51/+/FeT/
WrER07k7cc5oZMtyblNWrf6ONooYnlxcnSIN/jXdsr1QD0b3V6Lp3oPTLUqTi/xUbAgl5Pk1vEkv
Y408/8RmWxK4qfeiw8E5G8uBWVdu+ZcqaInzOcmVm6h6t5rP0uxCqwc/qSHFG63T0ZSr6q7VorcG
yup8RIm3K43ijYCBrVKmFoUGQddHaiaM/mMQqLtcFx6mBv7Y8SHVtAHY5MSIrCf0dCT/jMEfK1or
D6rQJk3T3cw8EoOkLKm2YZ24s6vp0qcoh7/71KEji498G+igLz6rg6NyZrDytOlBRtPE5y9tCex3
8QM1TjEwgW4HteCscVhTuHftnfMxOxMVZlYzdGsgG0WYiYtrIwdIxXaHGFNk7/gl9lLlhA3vIddm
QH1nSyvwAlCOoAwkqTPTGOGbWsOIpSLtVglHghm7s4L9hiUPDbCGO36FGKl0qpJk0HFmnzSeIJTN
7X61qbDHTo8G9ra0vNB7TcDI1Hof3ZuS7xzxvtcXMWw8xJtsEuyYh7WynaNilqay7RsEdWmC/H5L
nO2y2T2bd9m/32Son36mGx7mNAMcKFF8j543L6KR0B2n+4tStCf8sJhSmheSUvdnv4dL1VOd+ekK
W/yYhCXnqVm6fF9wQDZL/X1en//9ZxOQxSUtXmFFNXacfyqwnb73qiYiNBqHRQIHtG2muC/Nf+X2
vk1UakR+4KW/1+Sq/p6FyW75entVXmll76aABkDQ0tDERUaLNxSMDaIrX+5PLBN7svqntxR9ECfa
3WyavYLH2XQ+biSt0ReETOZ8MZi7Rsc3CqqlIbLhlAj0Zq/eoUz9mW0nzEeE+H2jzDUAVPvcwMcd
59bNewDyhGaPVSHDvM+SHtNKAW9LtVy84qO3g0uTB/FTqgZqND8DQ56rGgznwFXRkQfXRNUAmzLd
bByNw7Gs5dcO+XvJXrb4wBQBBahoX4KvB4ci6PfpiDB3qP9NtbKKC9R8CsfVsFZv+UeTcDKjOY8c
fkqjsNpWpAKNySv698GxCkOsCYoklKIQOipqltK6dG4/Upr812to1Os6Jo/hT43/C8XPj6NTw/76
NWgCLiQCOqKKV/cL6O3QttXtZ3JbH7tS0G4oa31buAo/6NpJ4zPv/1u778HDEekVANZKNbVDXHGv
BALEOKjmqO056SIswKy/tmL9M7obJ1NQCgK9gnZSckxWGz7T5wYNlzFFJ4Uiqy+zYDKbbDiijDxl
HMHLYolPYvLZ4dM0G04/sYVN17MY0yIFOTqp1QGIHAT4rLtujZs02KqEQOH4W+cGoW4+Y+XkDPKG
UIbCmLlhJ/mJWf5+LEM3Ci1SGFMygUghf9mqbw69gmo2cJNgj7EgvCL4O1m2fp8uSowjHFBQ7FF6
V9Ge6jezG0VEa6HHjq45k37z3fZLF7ZAJwloZR7m2lLeSJt3Sc4vyUxqagdd9g3pNY5iHTPVRuu7
y48Rb9+xEQkqMuwHZfAid0e6QCy76OFCfCjBIbEhRAETpaEukcnH6vAvrebTGIEkQHbpP5SBhHMI
UhtfnFvrHzosXoZ5dBo6QUXg5jq+0F2ttExiU6RSZSwoIYX/QGSM0aPsWkJGsdZoexxECkTm1bTj
qeP1//uk/FMO6YG+oWnKqbfAZfHSTKbEeGlN3aEfx1NZKNJLRhksn+Y6jiHdy5FU+N3uh1iKCRs9
ou8KYkIFItStiW1NkE9y4XRCY6Aa5sx5WGme4eS4wVBrGyjEglHO4U8wsbANvNKPNwv27BgBXjys
SoXsQnlGSMVVuF3H6Pm6wkvNlKJ3nwhdcKJpIBRI2wN+qMbB5U9dR9NtWI3s7wnQMlORDryFFBnB
3CyAyAjv46F6oCZcVpj5PmXkdhZnoIqov1Vb8L6LAWTHNNaCWRQn4kQIaSXkK8dzoedSf8vplpKy
QuRt3Uv108be870h2DbCFnmt+La/6K/B3u4AJcIGsGKMaecoHSfsSqi8yyRrKxcoO5nQCxYzCqRk
uIbETvYD4xfjJUV9RfGYcwUd7CA6soPy03uUwtDk6RvrhKWay/OayurxYscNBqQBpag4wtP6kGTn
W4IwFDIWM9ZwVqAvrRTWiE4Jo4xC7jJVKsGLtNK97G+4lMiVvTxLSxcIqisf4W9qivwi7xgAI304
w3osnrkwHUH/8rhPlhJt6p5BHGZZpFf95jG2El/ss/qmO6or9A9XXnPnmLxMlTQoasg+qZjWbEoR
6FkiXwHMzOSAsVJl7IhDNFbPvBVY8hVNA4h53B62taF6ClE75sEGh9lCSHozXrE0ZvKrxU2f1a3D
ahtqtCiT1lL764/oPgcX2M5g7TN5W7u6xzdzH79s2DqXeQ/lZYSs7F5oq8QP0XKtdVfUPDFcckw0
DTjdLGieCgeY85au0rYYa5XaiM0PXkOTtzwA2sXvCyILVsoeTFbBGzuwb/SgZl4Xlo469iP2yfUU
zCQDV/U+u8EUHpYFgsv7IbALr3cSgfAOYp2m/BLNL21snG5t/3wSQGqMtaUW3s9l09Md6PuDQV4j
Gc84q8Plhztfr/meK5ZZOidp03PQuadWEhT2KHL2kdunFHWDI3NRQMEvfqrGuezlEZQBNx3bkL7a
xRSyQPX0AvdtKWlrnZ3wgPhCJ3Sjfy9dJHf0vmJfeHCpRRf9WaCSJAW1/mB5hRpYwa28EcBc9z9D
GkT56gX+Bn65Rb6KAHYrTY7IQKI08auZUIdSCLnRFpkNm/eoBM9yIISH20/HzJKpws1dqzLcKOOA
271CJTAdFA3aoLET1bAeOCY+wO4tTPiVDDPB0SyrAby733uENxQKxbeAod9U3mm1aVBCLSpCXtak
/Z6LLDdrzRHUSHU/8K09DWy2Hlsb5i7x+jRbConkA2yS0BoP542vaulRYjuPQ5NDh4NQphcrildq
cl9HNEbeMs4yZ1lPz1qDESXP/lFHFAzczkaGT9hJBvuQ2hS3iALmADsR874pndIMhfW9lzcJGmGE
pokiMpKOTdunHPPwAwRj8jnOrtIzZxliTHvdo0cUdv7QJulVkC6BxHEFZiWui/95EjbzhUL2L/4a
SRNN3WJ56dcn7bOOc8pRZ58Z1DG3qj/FGOXFjq8FCwwFYqzSY6TVr0RRiays2lYqBgt9olCvVZ+W
JHcwTV+gViVeT5V97nn/SgWssgfrfqZaMyjPFas5QyjmXD4Xm6zBmm6tsPgLls9e97mtSn7QBJnL
AOBdg4qK7MSlN7rXDHudpX128ibuWKgwG/nvzGkpXC5TBrNSRPrUaxrYXG3zF3vaONGReHI0G1Ck
sXQ+oVJ7mT4JJb9228uq1sOFOXnOL/ZzNlI5k8TGsAzISk0jqGwR8Vama16wXq/Ldl4YwxwjSZJw
ODSCZys0plSFX06+9u9rhv5veIIG8Mpqozljjhovmw7kWtWzPKOT2n8B5sK9KtEfYoGalYJ7uRlM
3bzwPCPXVbmZ8iQvvtTaFm6jSaIFt1rCd6MqI0NhW/0eP8pLtcbhj3DEaTJhLUtvggwAVrC5bOT0
wd75qAqIViS+ShRiNL0NUq0Lp0RV91xnqdxfH0bhcbDrTjE+0sQ2qWfO4iYwJxIwJMwFzIMkfHna
8Vw8bCWDOoH2vXA6hrsJ7ZMGQ+OkZHsC/xOGkezqr5B9XHg/vPBB4q9re6pC2jonIJdFYq9hoRR8
hlFfLOYvysMnnqtTpzTuDHeGA63u5pbxvTlgtuPtaFu3LqaLE8+reB+VCGDhQuiR8f0vBEPqpkEl
3I6nAC5NnbMtD19LOomIFjjjG2LOBQNULtLXm4LVmTSWqcEgEbKHhKPR3+H7OKocCl7ZlAT31IbM
Vt0Zayv7CVXBk6VJ63jjxoXdcNYo1inzPzaJ1hEY/fqDT9V9Ue7x+Hv5vLZn8+TSYkkL79qsohag
fbpRFK1ShvmPRErGFxRHazIZJVHmQ3JeZnaotCCwAWXNWGDQ9E7ODho5yVUw0H5eDguGD9BoffO6
zmKO8UM+T9nXk6lrEcEanySBpRaR6ksIiSXrJb2G0hHguvSzQNYPKBwLlgJ8UGhTF2Smveq4k+8f
AnQVOAf1SVrKxQjNDEraFWihOyjMJhVy6mlgDpHigNuSvvsd6pJrA9avmx99/WtLwDG+G2sKAZ6q
ciLZTMy2o+iS45vhx+aHpgMY7X3JenhDBEK31uddXoTXRbcUaAhzhhGdUGoiPU+Vsg7M9yas5g+R
ZCD6zWeRunT4/sx7YwXqc+5o3dMWW6vvxOPcFuEa9+u1gVnMMeDV6xnqa0PboItBqBMOdTaRsvMV
vj792akWBEwZchhtg0BnOgETl89dhCBalXoVAqbqfRCHDMBhvcJYtns0UPeUViDnJdx/6m7Hd2Zo
Q79vRMXKWAJor9Jeoy07AUl5+ab0ZUyC6R0ROsReVYmUz+JcrJP8aRR2a4JMULLAvHyCbw+7Hgd+
Z8ECGswLWF+OjZ6vZVbuTx6YT6JY3XS/0fXeo0YBvEI/N4zIYP3D/w6tNa8qkSjC41LTCkzJwL0N
LIbTpfh8ACd6ThwalI+wKmz6YvQjn0wl4GilsrxKiq2xcWTc9+GsjZbF4JfZ229s7IozooMFP/Wq
b3yUp7xZwMi9lWa1G0FEiV1BCUxC4dJo0AgX6f0uMuuioHkC7ZscRVvVRdyJ8DfSOW84E6FmK+fs
rAMlyEYgLvya3oO/rqLfsDHHxZ/D0CTrHJB6Ix8YxS+BxOokdwyuG1lNuSSPECg+6Nhxw1HYdKMa
yqy9NcgLC9moVjAAzIj9WDUKjZC1NFnsKLIah3QsPHpbhmN/igrRdoE3FxjleqLxz+a/ZTN+mO7L
JXO1I88QQngIqOEaUvxo8HKKdpkKzxPFlkda61dZJegXZPyIqQTMuEgTuGUwmXwhCyI3maetuJ8L
KaRKtH9rxWq6USgzJFpsuL1O50BhQU6s+z5rrMCQ2EtmOnHeO4ahFCWKSDyakT3IZ4CyLg1TFmwm
UxdhWPbckT2GQiEht/p7OYSBY1elzFnLy5oNrSRQ9doao3NofNMBaYFkIdI9jk8tyVjz5xqRJXSf
9KAlNosrn5zNZtqvwJHJdWeD1UitSpqcu+OoM2RnnLqV4CQg5fUKoQ1XWP31GzPA35Y0/El/6vXA
h+LzVuZcsP/9BsQY3WVkNfUl+KSNKfw6PYYNE52aq8XWid3kq0fqJiXGShXnqzIwpGHwyZ566UgS
V6k+4fDoBGfROPqctRfZGPqY9m8JFb+oySF4swoBVbufsso/xR2hcgeUiljdzo7mmJRPrl1jyLya
kgFS88A4+ucw0qGriuh/NKjCHJqdOJO27xwkC1UpU2fGIwiJN4ur4SKDvYaPSAT8slDTFALzt/dq
IJ1GxYKebY4jFdMv0x4Ayx9lA76bTSUwO6Ktk7CQi0feNWb+Widf6NOpf87tuZH4Q6GnE7pFyfED
Hi/B6HZ/r4Jso0LqsTbWdmnvpv079Ag3FepdmcfbNQFrEBdOK9jqn8y4jrXK8qJrEzgqyXrO0RIE
Tg4NUgkXdORUwBOlXjXEUlv2LieBUOqGu4SELT6KojMysC03JZWuU5JLdt5OFJuqpyn/DmwG18NH
NY1Sh9pWbNIraU+1rix/SWGHzgkX4jQZwL60uoEfVR/xNJzRIENlXquVdHH0QmrpvgWJ4KH/KlWC
ubf4e3U9hPN2FQHhIhvALvPIwHDf4PstBuQyvnNk80SWQoYHGiLEYvjN2ArpoKr0wLiYWWEOOy2E
bbDYKNghhYXfxRuHsHQaDZuTMlcBYp1uF1Zq/xh32TPgF/B9L319nfOEXjU6YN29zPEXiqWB0s+M
KsAObDNkHu5RCuolKEHjFgjqbym0OVGEaE/fpephJMvoCQojx8v8iwXU7vI1BbS94C5bzgqf6WH7
5U07fWYUw4FVXZggwVA2Zzx2oW0udle6qB5swKFIoKDkasqNg7W3yrYBDn8l6xFCQ1iCARswT5EE
9Fg0DcCULLWjCoRe6T32YD6PlR1cGTOGYmjuWVXsWhE1dti1fmepX9YmxxsaZ6+fDDLNh2KqR491
xvyEEKPek4Q+OIKZmBJWFNnsVuSfSnrI3vwR2qdZ+ouCA4ZeaBVKm5U/PNBNfhmXzpJL3YV0KFFB
Y+46jcpJvpIwo8wa5xC1Vn/ogm7847W5Kd3/wIzjrwSHWsRwxd3R3pppmYLDyIBfgEp8fZcBw7Uc
g8pwSaGS+qTS0YVt7l6KZqTJanR/gKKzqFx0qfwS1doPjeQW0CKgZu0L0mCyFi51+M3s95SzgAbl
5iQS4t4zc7JXiJ+JHiMrdj/FZumjoIa4f2lDoaA8o2/fWXhU7kkauRrg/eSt0wn2gd7KwIUazNoB
XJjOBRl7uMFsm3hpdGjBRa1JzS8fxdlZvyQlqHlELhk7UiZwQAwahgNtM3Uvl4+pYSw6/ZlAX5VY
5DCylOyKz9ufYzEs69Kkc6RRPV+xVvb6wR3qz1kY86FB1dpfXf8vYN6dGv136WMStDtYE5jYN3Gp
FVdS7P2+Cn/bCd/d/AY4v8R7Si9YeltFvYbr1xlaNBMgjLR5FSQugaAf6Jh7uhGwhqEeOyytcbDS
QTt85rDRycvngIEIGnV+rzNnUAidKQXEOu3eQXem6u5NbvxVZrZEqq34M0xnJ9Hrm522P/nGc3Um
Hg3xdIP15YAdgv4vpqQPgcORSztO20jqtU5W8pvXk75VtFiFh5JfJVZb9b9xq1vd4aBUR2m5XYGd
FpSVNp8sfgag9Vf1FP2La6Qn1YjB5+zcd9dLO2iIHyoA2wNHYEIKacI3HkdLUJ/F8SbRoxeHZbSw
0+xkwRWC/eInV7ddoKt/2SBpYAG/7+FuV+8MH85pseHudQdXllrmF5EYZw01K5u13hoSe4OzCzSz
So+0H3C1tXoc25kItERFP36/NFvl2tYxuZ8xM3sfl7/KncNtgD8ovCgrQaM9hHOCODO84z4ECnWs
7htx4g4Jc2pVpfxvlltvFVhEDtR43F2Q24y52TumiaOtwFtA4QIyY67EXQP1ZgBjmadyhW7PMUbC
AojoX4yrd9OLOS6sPV19tAXTl7SYEd+dwO+JjvqGYJK3P4w0+ZJ9qncnjzD5NKZtxERAZr6jPuSh
YTebJVLuJBainXCVApCR+NrB0UEdwUo8D0HjR2iuOZgFY4HipYP1acQKgzImn2LCyu/tLr8EfCs0
/n+oBwb2xrY8gdaGlSsOGp49EfNL0//F7kEVs+gc14Ip7lf4FBfBHiwu4NWv3q9Oiwn0IFMuxIax
NQj+azRQXgVCqXeypwfIEJVv1JHnOJQPcUBOX7PLzdHHOG9JCUAcJVyFHF8KJFzk74onRTw3mmCV
2Q6ZazOr57F7dpj01xZE12GoT30TFjJhkx107alGPjyIVwFEi2nlYVF36cszaPqZhYFuWe23xpnP
JyUNFhKd/y3MculkixBoCzm8mX2j5G+AB7oq+Yead9HfmUxgx9qUp04ktXShvMgy+6HPQ141/+Hl
TTX//WhaF4c8l3Rb+G0ZsHzh+VYiBVdkxp38sNxS8KrK6CcwDohjNOawtBe17D/wlCVR2UOSl3AA
sOQPn2bs1hiifClNfkqmOifFWg7FzILELqtZ2Iva8ed+AXSeRZCECoh6/wa0HtHWzN2B0JNB9e7r
SC0Qwur/AZ0UiO2EQoQAhecEXdDzvPYKlN2B/5m8/2tb3H4VgFXz2gg0DBhsytKjxjRj7caM0FiA
WlutURW4DrTP1X5TAUbFzVQGDpJhx9fuhlOdFeb638jdRAPrq7PjVNuzNudUyaYCawHNf3PKUP6V
bCQfwwOaI3+EHGFqsh7IvQXLznxao/zOXNBKq6aNYTPGnhMmMaexwxqgbnjVH8ewM++KC8uVSLwD
8oZKKmGBFOzxl0zdN8+ul3bb/Vqaz3LHxP3LwTFJnk1iLKEB1IdcxdyEigw/q44ZE9DrtPK9R/4R
qd5cnxjTIVOY2eKCHidejqtBTyvKnHHmIiQ39ymE+39CeFVP4nSqXsnSgVNtza4FOWEUyrCL/yTm
N9AY0J1nDGnsXT3054kI5S2dv3BpDsGY2NOiqCkA73lQyFZzinzCX/A5TtNRbM1GoAM2wzgQa53M
c+HUiMpCMki5cTuagddzW2pkGFi+dDw0Fk+fmr0qJX4ASFMQu7BC1ANQ2EPam9d+Dkokih2dVUt0
lEOL2l+iXabJefHOQEG4IJeuHd3PGIbZ+AlYPYD+L89/iYpQYr1YXBimXST/vaTGusER1bc7Vlwh
mtBytp/fgPWE5JfuyXAcZiP88jf3OEIwZJ8vbI5QFP4RC8EAybri446km/U0tbWE3/b+jvdIgV0+
xfv1ILKUe2W4qZFJ3pYK+b2VyE/mKWdx68Cp4RrkhNrzpQ8V8izUsSt4/vP+A4xW7s07eDQUK8iS
dfSFdIJW2ZTh/TG3vfyjnOt//XxiJFl8T0njeo2uwql7ASvFADF2CMCHCNZoa9lrkND7TP9vlik9
N7T4qYiqDPD80qi6WZmfd9A6E5hDbVHZCdFpm31pG/h+66JyMfOJc0d4ZRJMDCuLImlBg8lZugvz
9zDvgYLBjtw0TahqMjA8uPCERwmHPnCNbaVf07ge8Px7gCNzqvnrWccK7BPocOfBJ+D391sQ8T5G
rqB/u1E9zQnOWf5jIELQ5aHOEKBp1kg40slw8OjY8hzB67d+4Fy7/kxOzE1edSYlkWyyjJy7ashK
5tqOhoRgfdVbMLWcgLxc2xEfhjSZjN8JT6QGJo17lZN8PSkJc/X4LhjUKpg0pRAMxXFAPNIspPBj
6JpTMsXxdCUCDlKQ3ipJGsgW71H/69zAGayXW1Iurk/+2PKT1Lfd86gT9jk+DyTOcSZrtNuvgxu9
L1Hu38MY1PS7ILfJBKajwzK8JTGuI2cdreEKKUF3HVaAa8treePxC+qht8cJjY65VF4nVGOnK/aF
IFoTZ41ZVw/M7tp2AC8GHSe2Cn2a5rX/1h4q+8Ako98NC4Zr/EnLYre1auzmkjsxa4qenbOjjrMd
SQ6hbR3qj30eeYtlhlAsP1514F3W1ePc55XhMK1stmSCJF8TKq7+QTVAsojJq44ipKZTjTcYY95Z
yRU3nQXk68aS6/K0qc1kcbVzmyh194RtPul6eM6YPioLeUDHc8LeC4M2uyIb+rzDW4IkjuQ6SQaO
KrU1yZyaGkwjeMIhKpbydNOD49eV3m84qMsnTEMUetrY8lvqTQPoF79qI0tsB1CNpL8egZ2YY2qf
zMSJ3XhBs4nrnqXAsTi70S8dFnl0X9fs0oNzDYcjE0rQxtplvkoDppccXFvQa+5II7Qz70OEWssa
ed4y3OVgroF/nJbZ+9GgH37Tz18hWJGh6PSBPIi512JyReuk2HB38sdoSRjakFgjtmz4eUm7tJ4E
wP9fTeqW7wfBa2LQdwaMPLjOu2wh1DUsUOfi7Oov1vvg8CI94NAe6VWN4JbiDef7MVIsd0WEWD/u
wh4CN1J2bTB63muEelsq88yCY7ZWJ/rDIHkIKqAGnP/6cAe8q7MfqbBCq08Q2XQDU5dryluuLoxm
18tsDl1d8xHIU7cmX+Xb8BxZJw/zRLxhsljUT9bFx5vJ4DGoLiwOfbZYnscgf/TE2on2KKhX8c9M
OF5p7b+2Urp1HN/kg+qlE23uBk/j6BEROmnlGSRUdFqdOtEhhUBxX8le6zf21Ep1kK+tryeNwE4S
pwto/DPhaLgpCj4OPWyXtnDu4kp93d/ocIRi+zOcDpstYeccjg9QJjbcetx6sLh2CGkFfPpVXiOp
xleo1TL320f4XTAW6lw/SkqSytfdZgQ+U9bI8JiUa5ONrlLEewatK+MJp/bRHTH63lTZMCyrN3bo
TAwYqykjFbF6PuBkiJgnGjQkZb8LXmsSUN1uhc1NlZqTJkuFJHUe62vAZ4Zi77t3tcrJYQ1BajhU
MJIaVIOoZVvS4QcXmRWGLVoKrqC38QRPjTIH7w9RUvUIPyev0+I2AVWhofgOsMVgKzS2DpJhCXHZ
XfFXfqIL/T64h2mTSlOV00lMHzgD987KMBvLOENoU1sumWnxVHkk166oxD8cSvj+NXXWo0NYdjMM
xT6+g0LCgsajDPKONDzXND+GPTnTqP/BymQJQB/3jbZFYvf1w/MtT1mqKpCVzh16naKS1ZmWpQld
zadrjr7Obk3b+FxjDMfQTX0M/JCjpuEK2bRDW/P3GAe5rV9OSQC1SVTVPDRB0gKtXnMTABiQAm2D
Jh2wbnWaxRfQvzwVAUkhpCqllyigtGrPxY4fhL4GrTXgO8DnOaSO5iWfv3PK+fXzkJC97/Sh44iQ
O1U8RLBW0e5rmdqPETavNzuHYW0TuSYREzgl08k0q7qjiEX6ZIkzFXoX0eyWXcMJvHcVoTwVb8XX
622qjzVDM12sd18dP3LC4qgrh8gdt4c8dktavqXnMyq8ja9odspTR0IRns0B7I2HeXRFJdk7Tft0
HqsKnap7Un0SoWClVBSM/4givpm6Ij9KaaHiPDx5/gROMEFOcC/gk3rOuYUdZLV4TFIIKQxm74tI
kqyUF1LMHjDYedp5vd0HgTDfJl1leMMHTdDhufh0N90TWIuWZ31wj7I2gcGQGLioOCFUw1znr+Bp
AV9OspLJ12kInrGsAVRqgjDi36iqluUxw94+7YuxEQoBJuJej2OWjD3ghh4LSzgJnzYjpo+I+1ym
CgHdFOETc/7RvLlBOhD1GxquyNEb5P0BdmZg4OdJMb2swFHCdQlx9dy/j31TZU5lVDYY3EiTmc6c
AWPg54pJBTZYu+QXJpOi8glDm8GcZM9x1hCvteOfXtYOqnjUCkN0XjD0mLnNiRAmxQG+BUTX3y3J
i5Q2WryzctkQolnsknE8uZ/KZMymrD622x8ru2JiXL861eMJPpbxOpQa6Kqk89HB9pdcv+jfvj0I
pGmf67amkxZwg3X3vkyLIOWyGVmrhShsavXnXjHNSzIT3exZVpggkUKUaKe8Q9k18ehgEwPYLLMR
o4jITu7NENdTBgK1KKnYVrcsHJ2rO2kUU/6YMStZZndN67Oil2LkQtzDMepriMx0Y/sTgJ6iJ8p7
Hg+NKco8NBcuA1dlYy5xI6FB6t8lTA8XkBEOtS3cegZ/F2wHXyfTRvOiaMyHsjjDclnxU0aGr6uC
YUkGsTZ2uIM3u0hJ4KEttGj7Q4WWe8YHCcgHnvkXpyBHB5TF9A2dw2rtBH1DKTySpqEl7tH34rXq
zJIR9MM2N5ZFDLWsEjJsJbvYwxbGZE/ttig4yNUIoLsZim0YHxIiMpbe2Kvmiqy9bUih3UMciDV/
bKUwmd3RI3HUmQnrxhWqU+p9d5XNzaaw7aL3ZqnYGzuTijHMKx77SkiwN1RkGZ9S1MxUfGuMosdz
lJ3icBJMdESAvCOhFayaG4TevnwKdk+F38LdoQDqZeZdAoRRtZzeVGgw5I17tViLpHBdQuqOWWYG
kf6/lbdZyICCeH5+x/ZPZ1R5NVBiLkBAScQ8EL92oPFGm2zj6+kfRDsys5UuoJfK6CH8NhHn8PJa
uF5sU2GMmBZ6dF9IpCSVD8JpylDUG232JQzbSXPGBPSXI0cvyAZTRPrAXFAKUm8WKKtw5FsrgjT8
zoBTZeKxIhLvwG/HDFg81hiw5gbSvsGHC2FWts1o6YgnfoG1kyGnQJA9NO4GPly+ss2egHYsHRYW
KkkBZdxc82kYtj2NY4oy26R3E5hlmj1EJi845W4v5xHkyw1sCLn2JFw3fQK1b9KMgH9FWavM4hyW
QukzksdyDjr57BiJ+6X25c+wRkDKxZgeFcD6mcBVk2e8kOYfEZGvBJmybRomZCdI2OOxVPzPEMK4
fedHVYjxKuN1vq8vjMKqeZs1fXv4loBy/vGAnMhaU+XHURPF5YixfnqGKd+W+T2Ixp4zWosETuRH
9M5pFu7WHvQx9zOpWGu2nn5obxeVhs50e6WuR+HRgKi297yfvLoQJ1GFlr79+ft3Gh/Avi3vW5qo
WyZXhbzD5TqSSxv5Xhw6ZOiHoCshZhVY06rTAkpTvsVJtf+diw8N7oHXwbL2Ml1n2OBBO/q/z7Vv
H+s+zsfdXOZ4p9JfDJjrBFgDSqTk0+ao0YksJzkPk3atR3W+i9P3Gu8/pZ1VD334aY+1MFC9BlB/
mUetgEmfdkaroSt4YwR8D/fn1R3C+xCwS0N/jz0zUqOStkaoMsotQ2BGqZlwB3r7yss+Olve93ec
/hscRB0T1JzQwFnQZo7c/bMxA57vZiO2UaBzC8/o/9kcm7Unofh6lZ1pIGyUnc/zTIUTilDaxJPh
KDP12aMsI5WNMcGYJ1VnQ2UJBEJwgSGnSS6lDwzXIu3gOtpNFO9EwDhzUhczAMXrdYQlNJW5+/X5
b4a8FBychzmAlFONB9e7WTARsC/GXc1XrX8ES6FUcxXMB4wgafccWjewJ31ac2VW17ps+LHGMS8a
5adcvyfkoSgEqYJ6DKOsZYik+NqnEyXphI8xj/kPeJJnOX/DebyfpFmfeurp8ULX8fsysQ6PwUbU
RAh85H0L75XEGEW5v60WrZaUfq9O9ypSOWtX5wcLZ0GwVUPZsklQ8HcxM599t1Xa55Klt8NCivnO
d0LKWjJlySRBkHhf5yHsqLGQia6TccrPS9BztTh8kUk2Ia41QXnkLrSmraaJnGlHt6dazpuFA9Gh
42Ka3OEb6DOnUZgIQaOUxR+ALUdCkMYy76ra7BAirKAdVgxitcabo4iQclKEc5hBmTucSe5wpAbW
o9H6d1vs7wOaHwGxkcL5989ChVmDgJGE5+PRIdoqvpTRsBLaZqkwLIIixVx80LuJDR+GSnlnmJ6T
7n3n4jau7+NB20N6mheiy3NUBH7ZBQ744G/C5JhLL36Y4TRyptfQT+lrBjfd58Ems8ylgMFqueKu
eWdFsDDAruaxGKdzPULdmiiqMdMsaQfywjDz1TR9JPlgUF7+h21+gKF0zDoI8cVcycnd+K5Ss0GE
O40x1f9xE2QGGLEaDjwkQz/sjT+EFQxZy8Uk30Aud70aFTaDFr8FXGCj/y5tKQL/G7RjYnzvWRjd
5c8i/CNGpe89y7hxCxrJd8gdpBMu9C4yoxka1Ddi8elSW5DA6YnOJv8zfpSJuOAIi9Ppz7Sikeim
OQAr+hdRXwdeMCHTAL/vxpyDARntX92+cNmgiqT6r/7FMpgVpC35fNg0uWMawuZQanbUjvSUC6PH
rQhlMF2AVgTmIv5yaiD+VR/OaRLjD6K6YqRecSCs1Yv0U4RIWBLWU2bxhOxSRVIk+fRuQwIG9Tfr
fVYQ1oXkaPfb/vafRFa2ykUSqYCfF9944lpq9jBTmXi02WflOC9Mm8oWDGplOulq84x8VLA+B/xd
4AKa2lpSelVjB6mnsoZtk42zmW3HT974E2jBFK2l8omjvjR2nk1VjgO/gfx0hemFAlibHtSyHgQI
O3Q4/z/1UV3iH2BMjIUDSc2g1hXBEJRZEI3wQljJBlr+ZhbCepdGhySbsyFBCsGnnGJmICl5KJg2
9zdaBrhO0fMFPe7bC3Hd8iEwZaeMv8UCYWpDWlEzxJEaNWRpjBVsiv4Jjp0oBhAMQsaJv+nCug4L
gBRVxYW4r30+w3uaM2fTqY3MKZ2uesxthybHRuZDmqRSY3drabACEFChyuP3U8RxUhmaKdslUW4S
O5VC8kAaSsUwWrHQ9G2FT9pLtF7Cf6z3t5tdXNlluJsEBy6FW1k8ON9ys90Ea5WSZR3eJop93Guw
D8h8Xiqm/FggYQ+ADyP9dQ4w0bsUQccjmGpYn2VJGlZGcLGMqP9pMhtszVok9ix3Hg++iZC5mdXv
+MsTZxsMThl29r817nSStJoeHdRl7crLxqSwsSNnJnNAV0siXU0HZPXu9J6GjRrNQp3BOU1qMBB7
omCyle71JUjwZhX57IQJlcmEzb0BucWTqOUw1Zs2uMFkmDGbeZw1Y+ABJpx/tkONuw973vCzfvzv
bkT9SAM+P2SDQIawIoZsfqI86pUO+w37eC2f6vaAiByEMIGnxYC7CptA85V34HemQDgbhu59apCA
rJuNV6bSJ4cl6t3aQTr5ZJ+XR8MNUE4b/ZjNCWZbqCkYHCjBX/GW1mflq6VzAYQt8/rqiIF2VPSZ
n4VTGTdDcNPcVLraji5566AlfWdXylqbJIiDS+ZFAtO/yhVN5MR260Tbxzw291cW6vl37APtOuAE
nZKWQnP7UBXyI+2CT3x9aIZOznGb+sb+NREc4iJ4fL2YtR8Utq/Kn5hGeXOFjn7Ncs4jw/OkCv8k
/SI+eiNaSvrSiZCuLWdgCX25QI79WZvBNe5yqCl9B7XVkcGA4px6GzOhEef3RRgceY7KTypnMT9M
V2/16bjFgT457vrBkJKip1zYieSYVMxSmjwVPFJKooqDpeS5licKmDBk6arSd/E/rZMaJvBYb8I4
qZAPEXeNo/iXAf+o25FQijgNCZd3/YtpdBkWJfTne1WkQAOoLV5HZgfOH3P4ocdNJbi/eJE+fQ2t
TYX614lTy9+3jtZVFIrifawn0bFZr2oG0RWpJrkitqKEvvKvesB3zs1rCDJjhkmBba+azO1Qp3bo
2SXRydfkLoDXo7LLA9gq5jMjULCqFm8QaAN50YBnPP3ZMEg8ZUsPCfoiS3kjuHRjSTbtLsHQmYYX
RJvutB9sPXJc/fTB0K9Pnmv6THzPWd9q4nQk7FUkof7MuaIrYYoXuFFoWNcEdrw0NMpszv9Ynmt8
OEgMZbj4HcKgPBVgezOES6kDwU6+ixJDOt2FhxzwOhG2H002OvHP8k6YQTcORnyr+PYnb/v0Y539
15sFStyMXSYsxNF/iSSkp69VlIEIYrGUpcmRu+BVH8dru5f1fYPtdY42b/GQF/91ivW1CAXVd2/8
gQShR/IV0wUayBpKXjmooxvrdRBnSa9pMT2xhxpSdEI4MlDy0aBbN7aAsoCFdDr2vu/LeCzEEIK3
u7hlVBEwcSGdhZQMFRaheUuT+5SS1pQKwFf+5AdUWlo5J83+wawl6t8H09ThtG5gRtKiA9Kb87E4
8TBV2OUX5t/15QAQbEdP9kPniU2FSZ0NNFih66ugh/5pjA0MT7M+qSSuAO+DLDHbEFXPhkPHqZYR
hQeEou74CC0Xo6ATC6QYWoFVZXKm2GjQvHqneVKLH1LVJxEwYoUkpqm/4mPmhm218Sj4hZ3HxMoT
qKjs0dQOI5M2gQhd2zbM1rzXPI5nzOc8iUvnHYV+0AMPxzFX26vNOKtIKqyuk7qKiKTuBTPaJXq5
mYG5pvqQMGms0cQQz+8O6rFpHrgWGI22kwTuI57MbK7hCw9qA6r6iuy5dSAmbG+narvnKn90pPJD
XGPHCz08Asm+tjJKir/rhxTabeewW5H4mulv0IskuzC33Y0rCNr1CLMqCjUXHfToEWsS6JEPkWS4
5G6f8RrZ8JiBk8Zo5vEGt4WLEDz/4A8qjMPnECuoQoqbepPLXOQAg3sz12g2JXLCvsFjqLBVvMYa
a+6t+kAYYBcChrRid4LR1DKeEYUsbrRAG0sxe3HbmsebewTl5RXaieXRl0bdFTKRDGeeXF0vU76s
ilKC56b5LpmxjPd51divM4pjdJI5fQxSFLE1cNqRWZnjVTz6CQSTIepPBmFOjUMi2iGJSxJEm6wW
8T0YbG2sUuaEf0yMKLZlm/mrN/RLumdkJZR/rm4vStfG4C2eaH5Ouq6fpKfYDyb3pGxCv01omNUf
gwvqgYh62/5RD9MrfoEhNfx00u2TrcOlzp4RLuOJ1EP8TWWqKD4nTw8Pq2bmpHO/IyfV25XeV45X
h9Nf4dtPm9wncBfk/uBEzOXZRA+LWjNuhI0Ax6FZ+6hJEAAal6ipxnJHwNPZ5gJ1s5ejHa9qSQEZ
Weg+TNdwGXxRvjmLDAL7MGj20YVnB3Kn5rkYDNnud17qAF8VD915USS/6fnRQuASKH4YPmCAgI6s
ysr1V+uXA5e8UIpK4MnYZ1WB4JwuTU3SmNa3PIXCmTul+mr0DW8/U5ELG0PVYFkRIQHDXvJk/IHb
Qwqt+HFfRhKtuqow6ciIIVjg4AjeYoEQQBkZO3Ua9+D71gx6n1mumZpvhWY3qU/wjoO3inXl6wvE
IyrtBfAChi4DgtujLeOX9fj4m2kejapgPzHKrcjj5jPLndddc9OvfPRlpcwug6il5TFQdTW7q5kX
0Cd6Z2eXtXTRbzTXIy9qKtV3QcWzALQHsCoXw1w7soDQcaXMEPAtQSEFYKvwj/GHEw+6lozcTeX1
bCH69U5tGiQ8j6390udB/BgcyrznQoOGZI5UPmhj1WvAZFGZVyOfxZJewUFa3O9ZBT5B9jsnAgtw
A55KwYBKZ7Am+/lYYqfAI/11J8R6cgQRKZLKICA0wLe94LFkABoek0HF5mt0rd0j5xkgVoYn5pE/
2qLANJ6jGxnJKfWpXIrGS5+n+CjsoI8L4bbXmwJXqwtu3PC6+k8kvbHB7Q5gNLgPR9vZhaShpZ4g
j06eKItvgeDf+LX2A86qh+co3ZUf1srbQVFt7uqMLDd4au53A+g4j955zQss5abvuL3p1VmjpMuh
3yEIMlokiHME9DB7pZrR9E6SNIwgAk8EdBpiPWgHpFg9ctyEcVyUDgtNpLdqyCYkFGc+fmaX2+Di
Qo7osCgk4eW/9NA6P8ADf2TA2LQCCDsvjTKwQMEBZT8h2gNJADcesHhRv+5MxEU8NGZD/+KbiHYs
xGwfA9wLLIekBybdfUMHI9YQfeCZW5svDczdo5Wr4NMmJ3JTy9g/U7nDpezUp/XLw41FQ+IaEule
jQOvGnkFqHTiZs4Lgypq0Xkip+EbgP9l5NsPIRijgSn4vZCHNSimYvOQM8TpNEbU+y/F5Fjlvdol
GharpUecjpPcKDwnxgXz1NY2QECTBLdgj6aNQOw9v59ntp7nlJK+C3x+eCniWvmLz1y6+bTW1NuN
kWDpazams3G2zQQZHW06XO4v5gd9TJl7+AhINdMBcnHrL/5HrVXce0y+Ma9ItnudmX5bh+OUc85X
JombOF6bBlZEIjOwOb0D6xN5UkuwpQFSoCTwnP+HWiSyFQJ76MfptdX4MxccdONgL/SNvNpYJb0o
rVax41y9WkQhXa11ULKFmSuLeePuTbo2bN+3hxuuBIAxP0gaesMtwedywy4sq41+VtZ+iVFfIRdJ
JUrH4c89zflYs+prBWt8BtJDrTKPlYAURRfA9aB7KNz0ZiP0wtyvGlLprXE3HWPe0PgsKYLVYhGB
AlW5vBjB90AM0rg+Lr0qdn7JUiXzgRCKWKgJ/yysavba+4jz3mYmqd4Qkby3ihvz86yCNFINpwYy
eVrVlVMzBfj/G5I5kjy8V/jAb4fiz6uqRVBm6NZECgDbrRlztMLCfMAVoV7ANfOyfzB+BmKND2KS
K+slkU8MAmIHYR5nAdAMKl5kuutCuakvQIS5mqxOLemQo+An7XusktKe/BxUpWVKcA9tM1foMYmY
2fRbQOPASBH6eVri7Tt0vtoEkpZt5TRUF1DBVPlFUFbZpPitIHCCXExSOMAq1sdHcAjC+27TGlaS
qJ8lG7jETjaC5xZnMronC3sZryxoNRPlDXEAmvT+h3rGace9Jx6SmXNwZKqWY+lZfgsKgfRu5UeK
kLak3oSIo/wMLjIlLKub7mkpMPvWcVn5+bOMlEKC+EzExaY/SBm78B4NhY2L46l2jAaW4sPgB5jh
sRMI0Kof3rB37K0xG7hRG9CmhLt7pDO8RUXRyOPjEGBEFbj40uccsIUSv52Hm9lVkX3TrFpWEuWo
MSw824w2pZJ36B+BzvNIt0x/Nnnf7lLTP82nr4bHZT9MzJmMvBojRAxKziSJsZ6BTuv4BhZuXyeR
cKSRTPSM0urCs20Ixzdi5P9hQoJQ/ymR7aBHmf58SMR9/sOTf7wQahRqMWt34WlwkG3u716MOWyj
RvbuB3Zg3a3RN4hXmKLwqseJE1Jkp2itN/Fave/xD28R/0/J/9zGbvakq2QTQ0jdAD9xir1uehW6
eV/M9zBb/TN1NA7Q+1E3MmtAGA3foUfErl8WcHvAUFOohEm1cFAcgxjXR6Ov8sMhNADB6Z639bCM
2LqSItvHSJ6CjSoWkOTwJE1LQUHBOlymkGpzQZRZZiu7G75lRMLeIj93a3gJQHR67nidw1XTtJq9
Nhh6MpA75mM83gTTK52WKalxgWWSHq4PEQrY2HG7aZHAciHrd6tL+SmX2Q7ck8zehTJs9URhP09Y
uk0vQul0brAGI75uNr/ulUqU40mnKqxExrjUiFfBP9cDnpwZSsweOxkv7NLNrlAErS3WnuuUSKVg
qvb99qz2Q/UKsFXoqP292Dybeqjd8aZyWjPBQOrBoEXi83s5x3f0+CbbAEXFEdkhrZxUigwmb05I
7k3NAek1jqT8K5xEFzMN0NsnPfbA2z68kW8t8C8GTjzVCegQh6xXOtfZzpLTn4ZvXgN9h7e8XbQ7
0+0hbGj9ZqaSgbi5pkVjtY6bsf82rJHlbV8oMwJm/o5VmyP2YUKZGM6XWDbzra6pV4hXAHiVjPxC
2d7l4aFKZE8RPZAwJtzOiC7p2onQjaCQ5/BO7eH7KT/kRT9uinsWfsq4lnAFuvBn0Z0GSQl6L6ne
eWjsUQumSsLU2fK+wQBAyrXshVyOG2EUEg34In0uhwSrugyHWil4Hl6qXbJHPgflb2Em+YkL695L
WjJbU1ufjwvwEjT/OrsAGs92sRGdXRX0MgNtBugJLk6o+EsLaZ8s+cpap4UONfmiEapDcQPpjSVc
SB2F8yiSepyCOr3y2IyN6zDGLfClJghZVjH/anBkDZrxrOpG7K4B3QLAhetPGLCqiiCFEFiQOCOs
unSDGuTJBle+NaZVl+lkGnZCCM6wsaQAoY4LYqd73hMSpx+LSn8uEtBJNPFozTujhtQF/PGQ8RBj
NmdQvE6SmPqPB0T4SCWvdOCrOStsphEGk6+ded1SmYsBOifEu2kywT+FOtfHXyL6ZUZoRDjeMll6
nc9NGfbtUrel+wKFENEeD7TM7SWVKjOvtbUPYSXhjkmlrKMsSrNAQim9rfyyM78eLzfuM083s07w
w+ytH5Zt5tFlxEQwtbYLrmi9vioWNmPE0O7k/FEpLyvYgg5uDIfqLubb6+vTGgzH4qCOgpZQBB8A
ckcoy8dfNy82HNdOgfkuI/1fudXbyyAkKqIxq9O77eXY8hl7Zqv2Pc+qyibj9bIAlaevzzB518ST
W7NLgk9PrM1wOWx8YDdpSnqqjXWFNylLxik5ZyzPio5X+zpVj74bnF9mblgZB2PIflioogSi/WIC
rbZx1c019PrW+n18XmUUb7u/xJwjQaHLFOeB+c6zxDqYE918aE/5BP+lqR39QdQo2LijfQH8rh22
6fe37s7/E9bEwC+09mTAdVkBX1N4iaT+eo4qieUNyaLKPVi/N7Fk1BRqLeRLUhg3CAbFqxDv0y1D
KHuI5ga4QIaCClIB2n6Xt+5CLLIw4Yis6en2kIGp4QV5GMHBYT9kAVEm+go0Ls7LUlDWbB/XndD5
zNaxLNGMg2mTKxHfwPUSmmZs3n0aU3eyusZAMEKGOdZ9Glu9IHljQThdGUy1rL8LfcZUd+ZCKbGq
bS/SQn/tkOYs4c4Tottsc8Mbgu6eUNgAvf64MyhuOZT9QKyJOl6b5ug9dIJMOhPEJjz46eejaa9t
2Cw9nTtJLdqk0pd0psHzLAIFOxBSsLWO++ShO35obUvIPOlZqDQoJs+Ws+hWCra3V46ZM0/ufMfF
4/sWbVI+PM5b9UdwVes+1tcKcdUq8Nl6yBSbiImDJhxQXNd0piu/boWsXmvm3McsJBGG0noCqQ3T
J+TEHj/rcMjq3VvayhO5dnXTsIEkRcwDJxAYrWduNw80QwOsPG0cmD2pWPKOQyE02OxnMdbA7lMW
wBnVG2RO34ORNJuZdPCHcPG8NVzSjS9hze6XWp1qPdx97BeXjJxMs9HjTsgb3NNOqdcCul1pzMgA
OKBIhm/ZKj40V2Pl3P/IHslKOeKC13SVap/lknKvM5z5UKr165BarwXTigvXKddyes/fq9+D9Vla
rUFp9OKr4F6aq2voZ8sOzmIOuO/IlawX8G7QBYuuz58jdV51gw+5Q7MLSi8Gzd0ct3fmwOxagrq4
KHBlHAn1Se6wjKcij90Efg63sgbf1fFWwhaQ/pT37kvUri4WuNVmlPOOxw9nquFXyvGfdhUu58Dx
vJlaOSa+rJA/POu37VlFMaKbq9eiW7Y1fxT5xhedfH4kXTtvPdoqpTIlY8VoupmeMHp2Q8Zn8M9F
Ra7oOOu2g4mwVOCowoGLGxjtNmLogBOXfNkUGrFV1zTH4E3OgxKpmJokRUCy1Id2YPJl2dH2TATn
r4JJdlIyS79yjYFAM7D7GjZTnBt2cepAC2V61BEHxrUdLyLaXY2nDJzrHvNmpUMKZiRfmXxa6lcW
OHdN4RjYM8lEUG4mja3abbx59maDc0+on2Jy1DwwvCHSZm0hePOQhttbA+YWLranZNhrs/Mg3xan
ChZPOTonTN/Sxn2UcbMrQhi1tWVCDmNwx5Z0cZ8Bxpa/AoUY+yYd57WCW9A/IDaES8ddLLFxXRmn
IHVTDaMIidNwu1ta5vhWS1xgUKif+83053clmJNs38/KgZicRYNFb62RqJEIUayzYHRDDaPbR8mK
neCQwSQJ/QBLkEmOMgxntWkx4+e11C7BQcLA8+0ZXSmHH7sEvMQqXzAh3Axcn3ejdXql1VptJB0r
W6C9IfR09Fi+BmlqW7Lq+wAo+7bRP8NMPPIJuUCPl7XfEApkh4uss+9A8l+BUb0BZs+jBbozMRJi
ijksLfk8Ane/s0a4ltxlGnQ6Jxn47fE3f6wLP/4x0JQ+Ivkqpya1BcSSgGS/40OeXYPAt5AVtqDh
lummPvFOmIEFYmDASMUZ89XQ+DyGtIGvct5//4/WN+xLctvxjs1BewfruKMququwYDGuTSPArGXf
t6jY8XgXYlnMd8v1ZL45pRFkAERZRcmqlT9s3FkGMruJlC7LmiaoEnRocEQEKco5uvpJ767zQPwk
9cBgxb/PD7Dm8QxpyPr3oTZko62qhSjaxbeaWSho3yNvQ1Vr858n4NjSOvBdED4AMBTqRM5EbPS7
t6rHyZAawbpTpal95XhQLu6xIXG2KgRw7OKF1/K9ZRbzi9GTYmSItVf28GHSBvNIIGOLqhN9enFA
biOHFYuq5cPo9Dmqt+R9p2acyfNU90gUUDM+dT6JRPP3CVGFJ11xQj5MCmi6mv17xvhAKPmwq9eE
IKWavvV9bgNJu6dUNo1fnYzAI927BUM84a2RTfdKk5+6ZjH+SDuaOHeX4DHxOoDk7oc+b3IHMj36
YYT52eIEzrwoFa88wJBMApJGO/71vszKO8LtSs3zewjnls+XwX6UXVJskZe2cr1NY6w79tBTpHWc
E4fI19ZzAeVkoLLUSS02FNOPjFxGS8sNu2KVxP6IKibFPlZ7a9S9gHYou10Svv8s7wEDqT3enq6h
22tAAh5YRE6HPamGX+/P2Jxc5H3T0Hzv5P5L7kSCCMctGhohJPaXU3Ve9GzspTE6UWQAnr0MRZO0
Bv5tmiumEQ0GwOEiSNb3n3wOq95Wmux13RJqu1Z32kbL985p0NUWLmXp15cjRW5fwfSf/E5HtiO7
imQ8cPyDTcIvy1HoXFP8u7qqvSn2Mo6X2P9IujEIrLsyQRa+OGND8W3zGtzd4mQhZyowvskuv5Nx
BaySTTa1tIPRpk3ESYiKf6j3yxAAetJEIbnoZChh2IofTAIhRVvj1UcCqtFeVZxbaXKTTrilyEgW
nSg6IsovxcJCh/S8GZpv63MKaOg6GbmJgNuZfXpBC+LK65Mhbbew/DIz9uNNeQkd0VY1Yp3OQIp2
qxrgioxE6BroQ88PCG2dDEAGuGwED9nJqgG6bROsACNN7tqCUX85+uY6I+B+a7LtOENmCvYD4n3N
koYIQl4RP+8gBDzchiyUAmoH0zer/LY2n114As+FCfCpm2m1DETX7h58JDhRS17EoBw/ezUV/XiV
7vnSLlWERRe95B9F5lrX7w6/JcHRSz0xf9E0q43zqP40PHgJ48UryeYqqMoD0JmIO6lFmBa8zkTB
qWLIHDXoi26LwlOQzRcLD/rYD7gR9i2w8xl3PyeeOivE2Il6ZZLNPm4Pal045ewrGbYUISZUAqk+
69KKUedoj52f3KQo0UJcGUnX2S6LAYSbvoUE4LS1MdF6YP+Vf+rYqm64IEhedo/IalsjcEmTrnQg
YOB4VoLQD0sf9MgHvpH/QEfdgDu7sKtcHdaQ4nnfzCRUkYzjleTj1MCR6qiCiv8ToQM+Isahm2BM
q9U1Ji8aqXoYnayh8fut/IJ66y/NcvRwqtkjgp62u4WXrVcnPAnneuLJ+vJ74o6EJViVtHRgb/FY
He83HtWNaJmrZO+kcdlx930tgDEpim1IIQW9bPf4Oe2L9YHc+9PsK3+ui5ve2QT6ADaAYHAKxvGh
0UwQmdrYgbYNGSerNJBXwaR0dLEvipBtqFRvsqGHWjlLcfm+bLdmAbVUQB8icR9FbwoOvwIFdbny
U/UI8lnWzqU2CsI+B/Ra/FkmohKtSib6xGVEKqMIKoVMeVH6LfeJY1gnhO95nUWoXVaDJmRuf/Of
c3Es6WcQaG3LcMOZsWHNpVd8YDuvcoJMfqH+1RLPrZCM2oEsRHYdCFKiG7vkAfRIvaQ10jjP59CR
fvwickhc3GQe9NBKvHSsBoUYHczwXGnC4Kmm0TsQQvgDa8MiAmrnTBKLPQYn1rC9/2eFmI2Prxjf
+cgBIoUVSyxtSjmzQRgOK58vRh7iulFyhHNc2JxP0lcTuH8jJjEXTRzFvx6lEFQ4CJOcvE3XIy5m
mig7yWDuB/u2VDeLsknpfMWq3CiODj5sNr53BEr3Ga9kzJem2iUU6DMzAnaKIB5MgjsUtOF6q6Bx
wXxSFWpTDQYTnT9ULPaF9iC1h8XP5tt5drWukPoJZrhMoKvklZx5dFQYEP6bgVMttIehJq7Bu6Eg
iPQBZSI9rCie/PBNZb35lk5wMD6ty8WEt4SaJcFLjPtC3fzOHtrUGZpfccPhlMSNOO3YaaRpuN+i
KKsET69rMB8DZZDIsgxbCvVf1ZdEY+KfCc4/plWmet6esSqZvQlVQyr4HYRK/XvSKZsuB1dr/dWV
Dwvm04+ujyKgv1U1HPKIBzLyWTn1npzYKYIgOTv7QbYqt4e7ibJ711PDAkhx8UcA5EdIqZcXJCu9
Qm6feTe6oFo0KtotMKPUlPNL3uBX5VuksGEDf2T2AdM7WEvO0sl36xM+YJF6ufb4SVO8QWfL9Apz
RWEmR8NRtAtfHrv1ut4kUTtiCf46acSnChwuFdyUQxPuVKuPbPxu587Lm2pWmMQYWBi8bUn/LHOJ
Xi/J/+O4oPMLrWjFIiy4q4paWtp9pul5amC+jqKEIb4KjSvt7KYlohKHJiZUVaIgGVv3FHT/JO8t
lFFa8D07vaptLqVlwfQR4MDdXq1XKQ5WSWdSmEuwZ6rgXeHtxltaTBsB55qOG9Js0m/vJHLMSAjB
RYV3VyWOlTnLSVcpcZ2jPvXo5dRi0FO+SgWaKaWixOeViaH28sGrFNp0EODNeDXY9MNHI3++ZjEr
NcpZid0UwIcNuTZNcRJeKNtwwQnl1jH24akAXZM9Wib/B9dWhQex8SP3LvhKCNqLqVCx0Hin08Ln
IUOU0nm22uhDiU7GcRxvCpvbMeNXY32V/wc5U0R6IFQhfF+DjGE8L1x5qnaVRYsL9FnPIDcWuuO2
pdrQbTQ5P1AHwOxdoisyd91r2nwAX3qKfGbu/Wr2p+a6CJQRTMF82RlwptvSK5+KP0sYQSCAWZci
6VhleJlSpV4UJGa+kGBr/NTAX/gRgJPfsLNqe34tGunV27g6cOWzTFi3ctybv+/avXxk6PkwNkZy
ueyScFXDztHs73amk2s1Lhzwq2oOY+oPHyMj74XtjmVoye3+acZfOGuxRdcW1wNGROavoQ2Vryqh
momRb43VTJbWt4inkojzUuxp6iTBHEHi+xK4bOUz//M5UuNbxU9n7lwkrrnyg/YVx3yFVZExaZHm
FHXyqaq2ePMXwnnZEQytjdo/8mW7quPb3O+ELJRAV0UQToQT7dQQvaZW0axV8UamWnuyAHRaNppJ
u56Y7oZ7ZjEahZ1+fH+Ax/LgF7s9WuNAAWZ1OyBwVLTCuf6h+yj3pnYWV0+OyCHuNeyxKsXimX2g
HQMK/RhYzJQm5n2U1zn3XPzjkVUrWP4gka2ql33Udz0i7n6mn8nBevbM3o2ElXLYArfhCEWmpp4C
U2FU/ClbO5hDto2IElVysPkNc1i43kZYxzM7a+Z1JUG4KBShQv31SXNqqDIIhyWIgA1QfS6MJcJF
t7Oxywzf1f2F46hhQMudeDmZ7Qvl0iC5FoH4bePtMbGOy1MPYbXxwjyHparRrmr1lX8w12WY5A1A
Q+q4stUVJLxIvmfhV/T1oVvN+LyGHfPWhkL/9oeYL2Vx3oj03uVvtF5C/sSrNuoLoq0BHFDvwH7X
D9j+abRubD8RJYJW6u3TVHtBG3ei/SG1jvV71XAiWnvT3CO/MET3tQbmAB02FFyRv6sPMBY/XJDu
Y8bQmZ30pDzgkC3qdAehssVc7mGW9BMn9mM7t1L66VcW59Vg2zvgQuJbsqly+zPBnkRSQptN9gEV
xfFikam5WjIkAyLUH6dKAQw6qw2CvRUlqFTEe3rw03pArld6Lxj6p8nZ+1dj3BT/8VZihc+Nt7zG
058ZFZb7EBOncaDXhLI9TPb1jHep4RNluAPZfZHHqqjl1BExzc/8l7LTcon6AHibg1Yx8goQpwfO
WVehaYwugMNDUsRp1YMDgK+jEQZTo5VCAbIWbb11OAE2M8aYVYiSkpe9e40ky+CmD7HF23+V7kFy
nmd8KkcbxWIg0262rbeeKSVjc5k8EvEQkZazspGw+zxb2lKm20lYdO2IqQyNGeZ1WAYY+TF6Fk+W
vZer7Ju2zo+MLaQ22p3swJ0pT9DWSyyc1vJHUsdVN27AhqjlXfGksHUJjoD8Kd674A36JDXjLP2I
yVtDiHazd0WbDy2/486Cwu2xruedg8KFKnIJp8EV1l0yr86N0UgBs1pHxr1w8LNiAQSJL+Jo/qNf
2sFVLMMFsktV2YPYIbJ1rclJuMnKnl1pkVL7EvfhvGAk3gkriTAXaV1XcolaHguUnCU3J7li+T61
1VSftxRS4ixUqNRWG7DOAHgqVVVSaMSfXmWQkRONpFAw1jPKdz/sREqpsKISHauEQoGymEOlwgxM
eZBrdHWQNlGo3NEKgSjU93CXf/sIZHwDuAIzSIUv8jiSGJ8ySvSb5HOanpZ93JMGQAHnlWS0at1Y
+wNVTS+t6V7NaFp1Y7JbKA3z2dmQ8VFPNKfNV10ODlN5iFqBubaK0l0lWHAAiUjeBCiMJ/2/ZBbv
sC0SbM/k5i2SlAACJBgxTAHXTE7Uu0tvts9v5X3sttPHbZBAGTRzGnYvM5nf7fuGVEPBbDtppwhP
uSzzxOV8GwQW5axmHEIn4/l17I3/DJ46Vc7fUe+jhBMVg9mx8p98k8XPW9enDWD3KVfeniwmxddP
AfnjbXXd+dN16GsjM/1GCDvTfm8V6x4ddmTWbnbjqmGkZ+wJ/xDz15SnSqU+x4F6Sh2m728uUL0z
40kOHcVPDJJQk8ai8ukhJSx8Lr9QDdQjTYchSRty0JGzh5T6G3Rovnb6BZUFzRxei9tcocLw4In+
lrP1t16A7TiexmglDn6kAOe1frqc8JBZ7AIxdPxZet+7OwC8ql8sl4SW7W+CZw/6Wueqk4e8a3Wy
wYJ/LMDeGamuKCW25jlZoAowxHqJ4Aytq51fxDHi+Q7t9x8KhyWUWvjDYntA4L34zE5XcSKnwaid
2reLRzWt4ZdsX0dU4/QDTfsOFndvKVHjatTwqdChRTV8qXVtwNBN7/CDbt/oaC0F2Lejkm4t/5yN
COv9RxlxY/WQdDelqMXL1G08NVDkqEZP1xiKa2VPpIStzZoiNKnSFCcq0lSwN/E4sqh79xYkkMSj
00vdMSPl6TZM+6SxYnVMzcWjep8Z4EaVYXYqC2fDGyK0QP23/fYtlZoL/hJakl8FZc7JGY2zi5h1
5QvniHT/e2vRfbTKpMm/a+OqHUZAWvVkvX4PoyPu3FY4tCbITwjLiG/yPrSKwm7pfJqUtyFzjM6A
p7PON2tt5PalIDeuTQhdylj5q8bJJCrnK3Mjdu+/nDDLOCA9blZ1K+tG22pdp0EdwFDiJ0/VbbTH
xEXWK6Y8aPjIKKMQZTOksjQhZ8Vd/WIVRapcnalagK65DDOzJvh+txFKpnSIGiBBPMUrPH7qOFPA
5coQxd9a+vsDlwCewa5ubzJWP1Qk/5QqbM3rMfWmQI1rOtVvb2IivTbtWwSkuA/VhnVz3ipvHghA
eTb3iKbsbfr/CTbrKSSoZCvhCJ/zOaY0G/cYfTysohtVMI92OtDT+OaP/Up2pm+IrFeG4sf7nKyx
mmpoKHt9up/jPFWTQdqGSBHZS7zN1dwsrNjyiFtR3sZdaCftPRdKoYvcYIzW4W3n11GwpiuVJdbH
SdskGIwBPiejHK36jYGsBtJHFHE/Ki0QVg2f8PCRAfKPlGo/YfqlZyFpSSPCJEiQEdXbytbvdJ7q
pNBY3yrVLhbuivkTLA87leNKTzBzjuEAckBAFOolKAcY3nFL7QHqWlMBhWsE4oG6LzxLuQyo2Zae
OZ0JHfWnUgZV1XAB0s4dc7n2HsD0rEFg3HkyWugJh67LXyG3J7YVvc93qBHyXaRlWyBfX0Dx/HXC
PezTH4Iwz1JvT5u1gxswTg3Z6dJpFVbp7r0qpqafrdhF9Trgr7P1bkaPWyCgRMpnepWaYSGG7Sdh
B4QHdFP2GVfsqnn0k7gt7nyUBzL22AMZbV05YgDIMMcPGSSBI1raPRpJnxAh9GYYPyz7SaWRIMYL
Renjggjm3Hz1QMdKi1veyFWUsO48TDinKii/DPqicevXQw8KZZhY9iKuiUh6VyuT2lGIemwVj1gL
18URmVVdj+gntUKu3vGG9mfT19dpowU8bleILSkm9EP9eWr4thxZQ4XUDIyTMXq+3k3gljkhbu8W
m3cRvmuN1gZ37R0I1+kebMoID8UrHVsUZgeE7YZsX/ZB+jtI8DvCLLyPCNOsm78/vQnq6i0pyVG7
lHsXhxMDPHd1o+5OZwC8wx2UT8LXMK5SW6PN5Q8RheCoHlL3n4TtKKUxUAEd7bXsdWolzrV+mp4N
z3Jg/5w0+VHUdqIExmYTiVrZ3mH0tiXcZFynoe6Y5FkMQSV1+jVhU+b1VsIf2Ch4hDoykpwWoEjr
XATwMdpVJijwIRXmKgj/FLsEC0He41HE8Nfr0IKc53sTMFfBTApHjRQeJoFiEzzPEBYTKtZa6k0f
aED9pxxAzK50dOSscltFM4As/qaigVBbf4LnRs//6S/92jRjp0x3yyZ9+FB47sF12hfbhlprTKwk
GywDpWE7y477SVHaaexzfhkPUf7nwmT7rhdU5fg9oW4yu4ZNkDjVwfXreNiFTQNai25V0Pu1X0sf
80BKItzoVZYTxIgChCqjgSfxbH11vwyibv8/7yIkIeM8XbALNUrIMnF4h3QUSs51H/v3O0n93wra
m7xqlznnvlWQ2zkk4CtUfG/G2QV5Om/GLdlM3UBZRUpuq0DZxSQnHlrN4Q5LNwMJkyivt8Lg6iQ7
O4OBdFUi/kMtrg6jYIq1No1g6ZEk3+HTzAkYPiWeT8ifUHqzYm+jaBNTmA8+Cqa+gEq5kdJY1TYX
avo4aU8q2ywccic+fm5Ug5dNeWLkLR9xs5g/Aplf6WDim40nH5EcPMN9cU3c6Q8Vpzlec9mhqWpR
8Zl3RQXkn5lwac4+U6h7VDJoHItaPIScKNnZu7tH6abggNqcuJPowgLYRAacIc0/veMVpcsC8eCG
g4NvTKnaKkEraa1wON9XusFp5okm0frtkMQSS3Jn6rwD/J30Pf6U7ICqwwHMRw7kOrjrLp9sDmxn
az68/N6dpPHm3vXFFvo28XnI8PmPq6Fw7tPAAQes+UZQs75w9YhrL4nFYjXsdzGQAWWyaW8cGDSV
j905kl5U2jBnz1dk0/OJC+Cq7SnI7/kv2ECnzny96Buys8lx98Hsu4y31drMtWuqbyCpMVYb7Z1g
MZJ9h2+3yOLJOGvyx65ZckJpUt74ZRNja2GzsNPIJhqDQzMFcctl9spQk3BkS343gqBlczXg2m3I
Zj2u9kxjGsMtZYG9Jhl5bR79A4vX+bup0GdPvUcrvQt6WXxL8qZHU932cLZcL1z/X1uZpg93E0K8
y/KL7OoQeBfanOXb0IGgqVRhKmWdMTCAsa6ESU3Wt+hTIvOdZ66l3V0EoLtiiNQmuclkE+FlCjy7
pj+rc8avQpbDuQpIHdGH2XvdZ1cTS7CZ9k/3X9hiUqcj6XPCQu7dwLzHGn2y/WDXO/DOU2LrKPiF
HDTdIqBdxAb0UV6bBOSwVvqzP/GYv1X+cddZO9/oVpA+caZMg+QiL0NXFe7xgKzVuuXwEZYFWZnm
1o2ctX1VbouFIA9Ba+FpPr2z9fCm3x3ermPfT6RtSNWahwvI/TZLpTYRdDBTGhJAIPH8tFdcKOkx
OqcvJtLPrIY9LuFCqBxhL6amOWDeQrTRZnssMXLBYYihdUu5CahJnpyaweRiMqZ3NkU0ELbUO5q3
yD9vWBIVtAznEfj6vrOOnTTiasJfNEza5Bc8bQ6Y3wUrPUTxM28ZmWbOCmGwso321MfZPAeg9e3z
QIovpSWulTeNmAwFNoVbXWJKj7siLT2SposjgKyILg0TsSnhjadyAn3RmdLDj/MdCwszWYx+sXtk
9x+ytVYtpJnCrx1ZZnwzHLfqktpND5h3coy7YVu8RlDXgiyDujzkB4FeLF+1szY2uRjsE80z29e5
28tboF8eITdtFcVuIKItwnRWCtOtOutvP7Yaghl3ArUbMEtwl2QSCh2dME5+YXSc2zlTHDkmHvpM
JiBdkjp2DbAzpDfdtyz5RGVDwGjp/KI2bIbd7v1fntXf6RF5OnehVskH8PTnZPD7/TL/5cj3dwh3
YtESvOTuBNDOegmbVE7T4hA1KkFnqYFA7rNWnLmBjdN2Nq+SPjpf5IB72jGPvl9WtzmKSSJ6mfcD
bVP+glAc9re2Y3T8Y63nbRrXAFoa1eywR/2HTwGH7rwVgmBUrr2fIFGRPDqu2NdlDelQpQfPQl6y
4oL7HylCSVy11BwW3vtfr5CS3yCRR7tGwIJIO7nkwfYglYvzemBfB6Wk88S+mH7Vs74b8d0aAPDX
P9UKUiVq/PebQyejf8qRa0xsg2OzGcDrnhJUO0/KMF6H+EjPwE0OE7LQHR/k0h6oD3NEmmWX8FGo
VqUzlwiItUva7o5U0ceejOEVg6WmV2JB0fq8DtlKZV+R16tp+MmoehwOLJ9976mNtkzgfMj6R6Pf
+BVoGrbq3GXswcSvAheylA+5r8zmVBTUfpqGzaNpTvG3oisLZ/hYQiKpmWlUBjEILa4PgfLHyxp7
wzaV6EuNIv+z5L0+E3RqA8BqNmJ/tB4TSqUomDaheMtid4pJZMr536hieBj3j0I/yoL6b/fQqA0I
BORoo9L0LboZqvYVnCHVavtcI8RAhcQg0aBVzOKZ63sf6vML1V6Dz7RhR5WrYigslgehlUDuVRn8
3pCJ4iDvLbwAlShRSzoyfHwYDwtxquDdf089NQh8ADdlcZm1SgB16HsUpAH14/qtScc4Srjszi6s
jtIY1Lr71xmxaM/OGbDLGutYEGpxoe9uV9vy5IivpXBfPwUZKfPZmx7x8Z0ZBkhApdVr9E05BSf8
w/lwA/FiGbpqdSjyhkCmO2azFTu/AU01HaGI3qcngWFQuKbW9ZLwnqiKrm/e45Zvnwr5WkuW9klj
dPlSlT+NuicKn0eIJHysHoXzHCqz3tNnM8YulOX0efemKudmb2AGS3R2s3bgLjycQNRi/Nep+O+P
IxR1tz/sByoZ6nmo9ydUdtPtW9ajkJ3TYxZwiXd5UEwSUbOKxrebCg//kNELGDzX2fXHEqLkDwS2
WY1TT19M5UAqg2Iwd/yGszg6+N8gPI6RlZ1yleoTkDe+zEN0NBHHyAn6BI4Q0tR2jaiFTMjq7Tqf
MI4ZZdNnEJBL3g3F1AtOLjMY1YBiWC7kkMpJy8weEvi5I2hdbwdwPkWMj/xHJd7l9BcJ05dUEVBC
vqbJH/4htQjBGvjGAGMJZMFe11gEdPjumw2u5Q2QGOO3Q5Qy673y1n0z4X4DqwmpP1N7cqeP1+9c
iRunI/1TR5gBlsWBsC+/A49FH8wpuflCh67/DwJqznUkBelBQqYIrZGZL2A1nnxJ65CdzJawx9Si
ImT16SZHjl+unCY9U8pZze+B0DeiHJdX2Z0dg8m+AkyaoVBlY/K28EB7s2Swje1/mG5sHkL9Sv3a
h+1oK/jQJb9fMUkAq4A1Cek/18ZmiT5p3PY4YWG7YTxkaMJQLIpOuIxXQxumz2erdJJ2JV21iMJo
54wPCN6BOvFq4Dxx7YEQnJyPADOEVl6zuCPe2StIOeFeSMTRgNIz9Fk77yoyg10QY5CMUL2L+hKY
V2HPzeZelkmja56Cp4upjgMDDDON9LSHXwyTvCrD+E9mX+zt+LnsYPHCjM2aTmbHFUIS2+tmopAP
Zv3mvbmfoTFcamtKJjGZFFW0eKn24E2SL7LzyynwrG57pd5FV4n66LWGvCSZg71+eQ38WEXp9Hhg
8rTZrF1icFR10OQUVyXR8VRVrOS/wrqELy8jeTqB58uyfgmt/1rT4l4se4V2huyjCzdEC7wenalY
AvVcrH0m6DL/lWw20I9nOxR1hMo7QdjSK9h2ZeiwcEUW6lM3d+aQNN+qCimiZGIFtfxcTvssmjTA
teK0qNPUmrJL79uqAAI1RXG7ZFcGF/GOcZaXvy4/wywfHxpmO2dahY/KAlP+ILm8VJPzxaHX90fc
vVwJt1HHLWuV978lVn0uIEb0v+b9s2XlagWSMz192sAHqaDe3mH1iufrKqc/4odZxkKLSqY36qen
w4oBTTrRdZIyk0LbZIEvQUG5BKA5NP4BuswVZP+l35nMy9ieJ6df/YWDWfdAyAz+Bi/7ikaPtyJf
PTcjRUrqYzIePVuMLII2GJ20duN6hzivWeXTMieXU1XfjHkG+8Lm8oeexvpIG71H3TcLJ8skK8sT
ql3nXFdRxk6VQl0gJFf4pOpRUKeuY5vsJm92xxZQVSE0qDCQsw9or5x6Mx9Hoy4qTgxSevmN3zzy
D7CQQTu+GYuDvFKkZgGMboKmrVZ4zYA3rqLyURkSx/8yZq6jsNQbaFjtrUkCR9feDduQaeU1aVop
owbIX38MNTF3pVPoY/FXn89ZpLWYgPK3YTimD1j7mOxobjhv60j7cwefy7rr+3lK3ESAWKXS8UZ8
6C0LRVcT7CLNBGinqs+KwJ/fnCdla7bB0vzlWzJEJwOwCFz2hUZcg6tUTH2lKJdSw+NdB+YTav9t
yFuMTDRtJkAYcV/+5zg0MAey7CjRjbRcODv6l+0ws1hCXqKA0/z9RTisjfvaMZCSlxhC458ThYd3
hJNHWevEkPbNjmkKzu+fvh81qKY3UsvIVhVdSTLlbosDVbt6iMQYR0E6Ry3wUfBbECh8AyQZhJ5I
jF4/EwR3j0QuL+7au65w4qti0oTlOApBl2ENMVVObxejUCbK2CNfK5J7tQsZPpbZ/3K/kYrDBk7z
BMIzpJHboJNbgWLiDgfAiKbnomqiNPSVFOqIba6UGBm2gL29m2oCyDVqqKGGV0DzwDLOh8o8Ni6r
anLIvhLMnd77coKJYb1uSG7CjPGUl2vABawvRT7FeUfpfazbjrt0H/qzNabw2/hxNg/yT/nKJErE
wMXbfhVOcEuaHSGvLYAk+iOKJKJwSbKS3We9SyBmeSsNEHu5hWqotsH4HrB/pHak3O7ai9raAkVr
57pcwTY3GH/fU5MhkdHpVM5Dh+Ez+wxmxm1wAQUbaYIB2xiDgPATQaGtJrgY4w3MJR52FNQsTOsN
6V7CvIuZxkN4KchDSbZ/1H3B3yDTEUxaoeEW+iTFWqor1ZpnymJy0qqFhAJ6QBN4aVMEONfwMLt3
sn26G9sv8bWZ91idxJ0hxBl2MNrruTX+gxBsGGfUclklyRij9tbHbW9fGNF4oeT3edKzc5mwDbjn
OvIzye042NrFo7DRmIs7VhpwXD/GZxmC3Tt9fBwMQFYkQNZ/3bbRK2oKAS023+b7vnELVJTcMDX3
pIdqKOY2nKbULaZzeAgqIXI4Vdew2nF69Ed0C15pOiFXFirEaTUnytva0kPlUeNlhVWzd7Jv5dZD
cnJhEt4I8fctGk1h9YpwfQniUEO4F6uKqv0ygss05wmRCT0lhAcKBx5CaxFPuU3iAJJfFqbqoyxV
QYCo1aEAJFRHv9fyKHnMuRFbgyh7cw+cx/78h2893UwTgQeyshvpzHvLCFj0MreXLLbncMDOU/mZ
J1axZeLYWvVV+vJ9AGwHabtgE4IJBfgH02DzrAVdpytZxrY6TjK0txflJoPkFAwBfmZHbWN+Er0L
L0z2x/ncJEf/kpyBK7Lp9o8j5BBzyQLbapv5PvbzcFYDwQLv9Rk3iYy6FFq5bPgNHUvrlzxWh14j
/h2ajdIuIeslORBS8kWI1aBzT36xZbEB1j5fE6qDANMN0LKE9vIiVRD4Pssx+9xTcTj+5VNg2g/F
iwX3A3VRg5J5KYZgv4ZihP0ExcMbjMO7QpwIrtfcHB9YnvhQF3NZQ38KsApbdfsTrS/HdwFWKM+1
dBCVZkwGxO4JfM66BDryFuo29CFAYxlQ+AwzzG0szWS8jutJcf/FsDowKo2Rr5AizkE3EJdtk3cu
3cmS46XbMGOinr+Q6qEFMQs3g7MX0Bt1Zb0ixB6Lk8jJj9+ZzfXkSSoGYgt2NGoV5/D9t7eWl1qd
ypzcLAfl1C/2OMswgAtKWPxtN5qCa8WYUgA0OOHeRMuhFRhV8bGlLUUQspv69zyh5JiWl182a1Ep
Lu2SFV6TXpveIp84fbWFB59UENtBnGDzQ7vcQayXt7MRxlkcef61HQhJsHasjsackyQV4ooF3lP8
bzKCxvk5H1s5EgBzGYsDEWpOF8sqnr7dIMNuZI0jD77tbva+cUfsD9DupTfSQLfqlN2VX36TIv8c
9cwSEMTedxFytNfA5Nyh47nTylmyO9tLZ0tib52KZNDBTNoV1nZP64znls8NF6QSbzEUi96CzRX+
ze/wYQnI3p3OZMqGAkRC0Mvc0IX7Wa5BwlQ0rrAYfQzn4AStHmsAg9s50GUy48MB39+F7NckEgLJ
wG03ek/qm0A9fF1llxynomwDzZE4V6xrBB+OF04yteYV/fG+8co5ku4iodg98BlfqMfn27UehIPZ
VRVvlNlyRwmH1ZzmrmhxB0Cn1tmohmkZse0nkyPTA+rO0xKzrbtLh8nWt0CTR+OlFDBr5n41KgZg
qiOWOTL2A3788Bb2Q4B3BACsErJMzd8VyCulk3JfeED2EAGCVw2jAiCL8ukS3E8UnhxKCmXczenv
b4D3lkxDW/2XvZ+nWjKoTFQq07ny3JyCKN6F5VfLrlut09ItJsFFtePXmNvmRxf38vetHeDVhSWa
PLHxgrgj9drEI669urr8z1L0YdYqHokPDtLtZlD4Z2C4nIrh0kybozzByJuvQT3HGdtBiLv6jnCh
dKqc5diq+qgHqZ67fGgN40pPRUZ+6wmRA6zM6i/XhPVobf+c5P65ZvYAKPJS4xp1mVbKxajYW5zT
KlEWDxe44p87tOh0L5Knhz1p93ufvhGmA6r+N9nhI6+qdIV04ukgXjAltfVvRvHZMNGh+HFGftRu
VvtrwGKDQBRNc50W0Ji3zPJZisUoA1mdbDcfNTw0JYYDL4/NRKjdlNK6wGxphH5oe+2HUwSB6SMf
v9Myi9iHMspceh0fSpzogPFLWAsUw1C7U9HTD+kqZgrd65im3zg65MhJUoNWXtxZEHSnMQtXQ4KO
TTwICKr2oGoHms95dhZeUCkhTfh7qLVw53otlffU/w1u9AYgcRE/1TC00qsW4jlJ0MbeVU/6LQsr
UIYJak0/kLCVJWDQ0gI3A9vXNJC5vVce89GXFW0kPMXkXnI76jM7H5tWi/NchudFFJE4392DXQvE
JrSAA28pkwEyJWgP+Y07uLFO0DM3IMFWLfTVglwOj10nWeviTx0tnUN7swHnhW9Rdko0n5D7UE4X
4csWTfbGOltaCcMFKIiKTFfMMHBsjiMLvC/NOb3Tc9y5yb/rV3MsZmgzfHE2ZQpQYCdC68xnyamH
XpPXW3ExI/4YZwJZDkJwVYyzdcltQ223+PUz2Nycnwk+z2eOZ43jwF8tjZcxSPUnQ57sYJfOQtB3
uDX2OyAG5yiB2wD51yRwkFHYqMWnBsEwK6CKTk3h7u8MwcA4X5xE/x3eyDx3XILK06B8+I++eSec
QITjh5ahcYYJeN3U8OwFsLLUiCKPQ9rEi5NetwC+pFMm2hCj+EOBJGYNpHrC5rNk5PBIGcFJL8bL
bx+dh9l0meAyqLog2TCDLeb83u4db9bh52QQ2jbXVV7UmmQV14vVvJX2Ta9ozjgmXb0DGk8Mjgsl
TUxMCRLNMzxBfMeSVmVEPvq6siSVtZLlP8qgJ9sOu6635MJv+tEE6gpFWdQ+p5gSoKIs1At8554s
pOvbxdkkybiLid6QpQdAFRHSTqmB+GBtcvegw5DnBB6a6eeGfCis+fH7ynl4njMQlp0YKuhw09Z2
HMYwHVhAdHhHGIrrij0+0q3/16PsduVO2m4FBXg5DIcYZQWwKJ3FABpXKbKzNM8OlNcv+ebXHEdv
iZ/6OujfWgM+rlJu/fPSuOGiQqy2/QD9SkKpiOzWqnP8P6WlX8IqdxGthh0lPBysNm1CegiLTm2a
cAIpYJ0+70QWXLjv9ekqDX5YuQDXWqFAr5aGDbgw3pnx53sGfjjbaEhC/elhmGSnr/wMO6Fi8hM8
3kWTjW2QAa80cqMxOqS4m4bcBIaVKmObG2l4X7RmytP4Cqr9ec9rFa7TsKsQTHZsYiRH7n+WfdGc
w2JMrHtCeisosWNwimhbksiHzsCO1L5NzI9iAIvoIjr8bfU2Kvt7ellVtrSA77FC/+xYbN1lKs/h
WNy3qdhV8B/WrujJUW4q3M3bSIWj6kRgIYRrxH4wDCpXUP5gIBJQSxMvaG/obDd8GHrNqdubO4FS
dSSbUA8/PydwodoXVKeh8+t+3h1tgAiqmAhIwnGs1bPPFOmmCs//aB9OWgH5jrXwtkPxQc0btI7h
HXk8swDQz1NgjWVtUNWSD5mPoz3m++kXp2F4hViss7tkEA443MNjXHOtaIiTzutETmtkq44RmrgZ
VgqaBH16fbW6mFvUFud15moL0VBpf4MCZBDLGaG0/X2WNmXNuvRinCJ12gURMzUu3GC7412HxMll
+g0iFgccXQJjPh7n6rUkS3FuTd7CucMm0Y8AZ1UMMahGB5ZH5JNcQf/IZGFLnNXtPxzYxybWs0g9
uQRf7mNXovZWIE8OWY0ipL7liweUuKURqfUZxwkGgm5wezqWuiAgbE4UyBUJsSCrmbi3b+CaETS8
oYxTAmQe4DPUlLT2lOMDK+uRjmpD3WjCp6Hb/ZbYSRSfOPVrITD1jZykAA7ecnEPWgDHkL8jMjGX
nD1MPYfIzRbb2Gq0jtGTSrD9Jja0sSqSLtgAjr0AE6Czx1zKhBwoyvTgz2j1LO1C28wVTsatXbJ3
J79NQaMpelQ2GwkZ/Ia9cfDWE98s7MfjYHd8Kkz8TxY/npQZmtB//GpkzkrAI0sHn3JcNipKeixO
yopVPw3z/RIMK0BAuW6W0C8Mr70yKFO+ws4SD3UN/1/seP7wpHnwKjeml8iQJxSLim3+zREa5PEG
NODDck0U7TEi1NvkxTrys/7jHa0GwSsw/SW0SpDOfU0WYoIWsNpVhAT6Ku2JTvRONCAyBvien9L8
FLUUn/R6dM0ptP2VXCpyRCdO5mLgxcBPNAtIJpKKX6hOQrhgzH1kZnhnRVbuFYCXDJmPS5tdRTC9
2VGepS8SfNYhyFe5r3kl8PMt1+Nkb+lwtHdORBLy+/ItkgWxri+0GQH+bheSgdN9PLt+Eqze4sis
gn3Ns+GgwKiAAlGBKoD2K+s8fZcrG+9eT0h2R4iUOtsfaFk1sSgciHdYEr24lvxLUdG/5OZK/UdE
JOcXhazbxa/Por/L1e8VNfdynidKVletsnGgldKQedWPWJ4KC0p2Gw9V+qZkerQbYfdETZKpHbVs
nhp4YHVW1RSp983IeBaKa/bfEC15gD3D9PumHT6UwKXkAkWIX6r6/RBiSPpKKCPoqJQ+IEMBaoNJ
RhUETsCj5ORS4GWcdbeMylDGxT+soM796OqPfJA8Gba+I3JjjpT6yFk5MU1OMmXBEDvswlQzRRJ4
PWNm/cBKbdIAPMnbInOhAqByqDVCtY9e8QBEBVj2n79HqiAytEq/hmDakS+ki4fhpK01d1ua79rN
VJmzUaa1Rog1b7chmSasqnp7wZsrA1OmtTWBBjmaO+5vowhddUtUm16xq0WY70fORHAJB1SWAsiE
HHZX3vSl/zFJg2A3LJw/OoxgPKA/Ta2Ya8erx9q4TfTwyzwS59z8jxp2d5itPf11zBLyvhYEK2uL
SOi45iEnQCPqtmwCOYc/BR1c6QOpYXMfle1q7El4fnBR7M/WmD2Z+kCE8GnBDtuUmMXyqp1LWXYZ
OB2FmPvV1YvVrEarKS/rYb3+kJTwZNbUznjM0cjRfsuXH/TejEiwzypPfx9qif6ciUOz43EIylcR
esBVAK6H33LSa4h9xiuPp2S+YGJrNCef7U2IAGTNcnSUHVTdSzBQ6MazIjYCmAaql3S5+W1LmlZb
e3S+PADL76BZM5GiOFGaY1PuQxogbCGlJ33++iSZ4AQnnM5xSSSE/gxIXIdRWXdKPba4VDuefy4b
IA3mBBr+7J1tqZYDzIhMmK/UFXeNgKCL6uDDW/tqM6QOzPM7mbNl7XZ34LH0xLaMLg6IIyJm46Lb
s7MfKC96ahOB0ZImIe/RtGaQ01Ghk2hMBI1tHcGlYBthYa6UUghAj8J3Z7dpDm3Gv8ZDhDU3Bseq
DotAzgkqgDwKKSV+IKlKPPRXSE0Dw9lr65kT9xvC6PWKKr4zFe+Qvzh/WbPQe91qyZVL2mMVm0O2
WD2EqvYQIddUTydFPMiNGVxfVgbio/zNM/o6QJip6Ao4GoZ0xdq3W1smDHItB2rTY5p/TSHLa1M+
1qY0iKYJSReYtdECKgQRtObJBiZbbpoEBrm8UuLYkDPN4AleV1OFYPGCFP9XnfhJMZGt2gkzaLZ+
M/i8jyW8UXJa5ETSEClMSRf6Ej2uHmEsFV5+AbYyxAKbtlNsBBvRa4BLCXLpmeNpubDJb1135mwt
GoECr0UoUUA+vvJesYC/tz36utvQ3pQ3wGM4hls/yhqOMXRZs6Qzx50SEdpgjADLEDUxezRVOTAQ
r3IX6N4nH6mJzbmT4EYFGoxu3RIX4u486vryjbqPdAr8+GKdUyAj5CiOWLmtToPtErTnQxEeogmi
0qdVhXi8qN7An7W5doOedTvCy6SG4Y4daydiHX+H397sEIGZhz0sEuFS0eQhwBDhFDvhpwB1t6G8
tlpkqrDzgGi77UxjXP/JhbdeGuceUBNzPkl0U/Q8Cxx5zrWEA52rMOqYePu6pb633yP3ai790Jni
a0npx/43Nec1WxiFHdQqWOamh11cODwGuDiAGh838QjGr/BGiXnB624yh/t4sIYaK+Ab6/wciQQN
93+fgPugR5RJQG3CDmoVg8vb4JkSLb9Bl1eLxQzd7VCZjwbbXnijaEWKYVkuUyBfh6eTQhx5wsDd
IhC7wTfOkEiuKlmYtmxCmVbVvqnZGyEanH2Oue1O/0K+uIcxOHFzq4WhOomqtOsUGNWc7a9I+cs/
VHNzSJg8RItS6UCN6GysndYjONJJ5b1T45Sh+cli8WGvYhDErgKRsAKGVosFVgmQZrH1Pn6skRg/
RuOOznoc4J8x3q3284F5SpVHUMSXXjhjcdYWMF7Xy1QnP8OwBP2q/SkzZH5Vn3XOGbIHf1l8Vmhw
ifIasbMN+lYE7sj9/GZYZqORTLFD3WkbXgeSWXs5cGprzyjDs0LEWISMcnlb+EfYd3xrtVdTrcYd
Zmw381ZSOu0lf27732SqtwJI9l3YDDecRJ+zgt/krjihUi99m9F3cBALueKd8ep8nhAur/AiAcZn
NBDak7+dQV8Hi4hekfDAKmanXY4mAVW269sdoAI0Y0f+OLD/Ls2+K0LF+vZBPYeTggS0wpjVIXew
mqNbwIKACdAMzvKgxaO558rdf5jrC5QCFjBBEJtXCT/V6b6j/R+395RKaluqcDca9VCU7tKozcr8
OP8sGLTj56S1OU/Q/eQ8vN4roeqMueQtRFPe/q7yqAWVyETrxDH1ICC+dQ2mKDO7P9FPm0golN0F
NQfvbkKe0at5yUF4unF+yo5J0TKD0dOq+ap5e8ZdDXxzmcyO9ywZW1DXsPgQrHPRHPnkb00Pz2LF
IAQ2CWvjYKMZaijEvrkwfQYprnSRzTMAUxmuOdGjB1szewhoDdz0LFLqLwJNOecHj/1z/EgcYee4
UqdTXc3KgUrLQ91JWyEPWrxWqyOm90eB1Tq8lU3QWioltkEKDeFfyTYmTTMTO4Kn29T5o+ZVZIrn
TihvHUe9XhuU9a2Wu91B4zi8P1FUzP+wfhec7Am5tv+MYlHf4NYvEbwLJjK4pZLwKg6g/spwAAgR
MeyxqILYRBNflDsLElgeEyMNuxI7jL+NtyxHCgU8hsy5mXCC/j5RXvROr/FpandWVM5U2T15bLKb
Xn1pDgVIcfblS9cxHey1rikR3rW9DhkBCK4+gXFOGCzR0FV5WJFvkHudGpkbSjWXTgQ1PHR9OHRo
O2KmEH479T4hURJ4pjueUlgO9kRenpVEOZpiwkr6mmQoDumu5Y2CFNOJ3heAx3BkBaFa3hZNuBDl
orB9i8YHQ/fxD8ObYHA5tz0LQ+F28UqlZT8fi06ivy63wdEdHrVyxS9opnCMPM7sDj3xLcvdonVL
b4nczfHmxi0p42Z1/Bp2DMsDdPW1lHykz61spLanZyC8cp4imHC5cZciPaFcnNWADKx6R58xxUxy
m14j3ZtW5LVPg75R0Lfexeyyu/2v811ePS1CgCWNlRbjP84TBYRGs1d/Hyux+z3vGwrn2OY4ihrh
Zdk1+KAVbt1MRsnugN1Kwc9zxHGfzsGQgN9/iQoqkmgV9iZL5dtgBgVd3eFlJ++vKYHYeqxDagst
CGddsAIVzTB76x4P35ABXLaBLsas8CdVOjrmEO2b2OrN1Xdeu1U8g6WLPkzSsayRqA598CG3CrGY
c1eIy6nhG57xLyneZHpcNf5/CAO0OFeJzrEOj+4e2CPpYAwVq1YHUHqQWP+cYOHzFHGvQ5ab9GNZ
HpfY5u7LjtMwlo9TGdLtkBfGj78zln0PM05mYUwUrNC9rBJzu6BX1nluWfe1Ez9ggfSd/5qrbeEv
kddZCDwCpMDK8PZUpwmirqDD0MaPaUpRqRxXBMizwy172pyxegAQrbi5iHsUzU9R6htqF5qrD2dP
Vlbe+HACn1JW+mZSsLbbIfnvqikV6z6bJ3pD5QBYeF/+0BeOXI6JUwzedHHOQSBOvXbGNpBIL0iM
b1az57w9OCRBCDTfJxZrheA/If02vGYyc7gPtOYMvxHZpY8Cv9onF8DLfMvh7/+lVX7C7H6RWzV/
2lezSwBhQKF1ZECJs6P4ardDVzV/jGLrBuZRpQkcaGzT1SDFLR7AlMK9maqHRw1ebUOnK2pdkTPF
dm7vb0qcg9HrnQqKJkNuLc/3KMIzbAaxcTgn7pmxGHjugawlRnLb7mdwZ8HeWwe6PiyUnMAnxvL9
oIraLJ2sUv0mTbx4Qyy6gRt1kH9KJlfmnTERrpC20S5WOrtSq+pszx8gJsrk/nd/2w0VZ28Obch1
RR/UJEtcV77J3A1b6cIP993bv6Nk1vYzNaApG9V3ZSzai6vWq45duO2nX+KS+3NRZcNic/OHYtcE
0N1ihQ0nCMpm8s0rXpynA+ZKp5nGUUMYF588jgFyizx5OcpdNTjr606Ws/Y+jqOP3E+PyhkpWokK
dgTXq4o1Ub/VIotuxgEyhQp46n+MA+m/Dvq/D2VT6x9ZJKTchYGXrYKd5FsENwSOkuX5gBLWl3Ld
BcNPf0dDnZvlpsiGlwQto1u/FOO1ortkdginnnxUIHt2SZIoPQl8A4zcplazADEenC3CpLh+GhWt
KQ1tMy7mIFIeJjmdI0X2IG3sngiWDfwdDAdHPl9fgFl7WOKvigW0s+7SSohTDBzvQzH2YQjOD9Zf
W9bow2vdNXhWTKr5TsjIxhyvr4tnC63iT/gYaNbyrr5BU+8xwzkoAWxu0eXbFE8JDKe+uGrxk09H
/5mADbKap9WO25hQjiRveuPu+Hc9E8Zt6xWftFaDFXCZ5L7ZJ8zPL+ujXJ4nkAG8Uo9EjJkAlRpb
0Q5sJJNi8n4CQ6xla+B7qhUA+2BZ9/2/zEtouNRfmElFIeQmOoCk2oSTObmNRZJ47wOaUN+txv4Q
7+tV65aKEEs+vcWZfjMhn+Z8tRYIKL1rG62YQHMYCFqByXqkrHY3h6dcwmBRD+xCE4ham0BGann+
fEpsdrarbH+B0aTcAnzoX4XgbHVbYfJ2uFs7K6Swk1f7aD5RviFQn/AWCf3sdKTbXBsdLyRvOode
Dl+W4jsb2MLSyHP47TDvW7v6aRt3JG+u7ASelAY=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw5a;
use gw5a.components.all;

entity FP_Add_Sub_Top is
port(
  clk :  in std_logic;
  rstn :  in std_logic;
  op :  in std_logic;
  data_a :  in std_logic_vector(31 downto 0);
  data_b :  in std_logic_vector(31 downto 0);
  result :  out std_logic_vector(31 downto 0));
end FP_Add_Sub_Top;
architecture beh of FP_Add_Sub_Top is
  signal clk_d : std_logic ;
  signal rstn_d : std_logic ;
  signal op_d : std_logic ;
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal data_a_d : std_logic_vector(31 downto 0);
  signal data_b_d : std_logic_vector(31 downto 0);
  signal result_d : std_logic_vector(31 downto 0);
component \(FP_Add_Sub)/(FP_Add_Sub_Top)\
port(
  clk_d: in std_logic;
  VCC_0: in std_logic;
  GND_0: in std_logic;
  op_d: in std_logic;
  rstn_d: in std_logic;
  data_a_d : in std_logic_vector(31 downto 0);
  data_b_d : in std_logic_vector(31 downto 0);
  result_d : out std_logic_vector(31 downto 0));
end component;
begin
clk_ibuf: IBUF
port map (
  O => clk_d,
  I => clk);
rstn_ibuf: IBUF
port map (
  O => rstn_d,
  I => rstn);
op_ibuf: IBUF
port map (
  O => op_d,
  I => op);
data_a_0_ibuf: IBUF
port map (
  O => data_a_d(0),
  I => data_a(0));
data_a_1_ibuf: IBUF
port map (
  O => data_a_d(1),
  I => data_a(1));
data_a_2_ibuf: IBUF
port map (
  O => data_a_d(2),
  I => data_a(2));
data_a_3_ibuf: IBUF
port map (
  O => data_a_d(3),
  I => data_a(3));
data_a_4_ibuf: IBUF
port map (
  O => data_a_d(4),
  I => data_a(4));
data_a_5_ibuf: IBUF
port map (
  O => data_a_d(5),
  I => data_a(5));
data_a_6_ibuf: IBUF
port map (
  O => data_a_d(6),
  I => data_a(6));
data_a_7_ibuf: IBUF
port map (
  O => data_a_d(7),
  I => data_a(7));
data_a_8_ibuf: IBUF
port map (
  O => data_a_d(8),
  I => data_a(8));
data_a_9_ibuf: IBUF
port map (
  O => data_a_d(9),
  I => data_a(9));
data_a_10_ibuf: IBUF
port map (
  O => data_a_d(10),
  I => data_a(10));
data_a_11_ibuf: IBUF
port map (
  O => data_a_d(11),
  I => data_a(11));
data_a_12_ibuf: IBUF
port map (
  O => data_a_d(12),
  I => data_a(12));
data_a_13_ibuf: IBUF
port map (
  O => data_a_d(13),
  I => data_a(13));
data_a_14_ibuf: IBUF
port map (
  O => data_a_d(14),
  I => data_a(14));
data_a_15_ibuf: IBUF
port map (
  O => data_a_d(15),
  I => data_a(15));
data_a_16_ibuf: IBUF
port map (
  O => data_a_d(16),
  I => data_a(16));
data_a_17_ibuf: IBUF
port map (
  O => data_a_d(17),
  I => data_a(17));
data_a_18_ibuf: IBUF
port map (
  O => data_a_d(18),
  I => data_a(18));
data_a_19_ibuf: IBUF
port map (
  O => data_a_d(19),
  I => data_a(19));
data_a_20_ibuf: IBUF
port map (
  O => data_a_d(20),
  I => data_a(20));
data_a_21_ibuf: IBUF
port map (
  O => data_a_d(21),
  I => data_a(21));
data_a_22_ibuf: IBUF
port map (
  O => data_a_d(22),
  I => data_a(22));
data_a_23_ibuf: IBUF
port map (
  O => data_a_d(23),
  I => data_a(23));
data_a_24_ibuf: IBUF
port map (
  O => data_a_d(24),
  I => data_a(24));
data_a_25_ibuf: IBUF
port map (
  O => data_a_d(25),
  I => data_a(25));
data_a_26_ibuf: IBUF
port map (
  O => data_a_d(26),
  I => data_a(26));
data_a_27_ibuf: IBUF
port map (
  O => data_a_d(27),
  I => data_a(27));
data_a_28_ibuf: IBUF
port map (
  O => data_a_d(28),
  I => data_a(28));
data_a_29_ibuf: IBUF
port map (
  O => data_a_d(29),
  I => data_a(29));
data_a_30_ibuf: IBUF
port map (
  O => data_a_d(30),
  I => data_a(30));
data_a_31_ibuf: IBUF
port map (
  O => data_a_d(31),
  I => data_a(31));
data_b_0_ibuf: IBUF
port map (
  O => data_b_d(0),
  I => data_b(0));
data_b_1_ibuf: IBUF
port map (
  O => data_b_d(1),
  I => data_b(1));
data_b_2_ibuf: IBUF
port map (
  O => data_b_d(2),
  I => data_b(2));
data_b_3_ibuf: IBUF
port map (
  O => data_b_d(3),
  I => data_b(3));
data_b_4_ibuf: IBUF
port map (
  O => data_b_d(4),
  I => data_b(4));
data_b_5_ibuf: IBUF
port map (
  O => data_b_d(5),
  I => data_b(5));
data_b_6_ibuf: IBUF
port map (
  O => data_b_d(6),
  I => data_b(6));
data_b_7_ibuf: IBUF
port map (
  O => data_b_d(7),
  I => data_b(7));
data_b_8_ibuf: IBUF
port map (
  O => data_b_d(8),
  I => data_b(8));
data_b_9_ibuf: IBUF
port map (
  O => data_b_d(9),
  I => data_b(9));
data_b_10_ibuf: IBUF
port map (
  O => data_b_d(10),
  I => data_b(10));
data_b_11_ibuf: IBUF
port map (
  O => data_b_d(11),
  I => data_b(11));
data_b_12_ibuf: IBUF
port map (
  O => data_b_d(12),
  I => data_b(12));
data_b_13_ibuf: IBUF
port map (
  O => data_b_d(13),
  I => data_b(13));
data_b_14_ibuf: IBUF
port map (
  O => data_b_d(14),
  I => data_b(14));
data_b_15_ibuf: IBUF
port map (
  O => data_b_d(15),
  I => data_b(15));
data_b_16_ibuf: IBUF
port map (
  O => data_b_d(16),
  I => data_b(16));
data_b_17_ibuf: IBUF
port map (
  O => data_b_d(17),
  I => data_b(17));
data_b_18_ibuf: IBUF
port map (
  O => data_b_d(18),
  I => data_b(18));
data_b_19_ibuf: IBUF
port map (
  O => data_b_d(19),
  I => data_b(19));
data_b_20_ibuf: IBUF
port map (
  O => data_b_d(20),
  I => data_b(20));
data_b_21_ibuf: IBUF
port map (
  O => data_b_d(21),
  I => data_b(21));
data_b_22_ibuf: IBUF
port map (
  O => data_b_d(22),
  I => data_b(22));
data_b_23_ibuf: IBUF
port map (
  O => data_b_d(23),
  I => data_b(23));
data_b_24_ibuf: IBUF
port map (
  O => data_b_d(24),
  I => data_b(24));
data_b_25_ibuf: IBUF
port map (
  O => data_b_d(25),
  I => data_b(25));
data_b_26_ibuf: IBUF
port map (
  O => data_b_d(26),
  I => data_b(26));
data_b_27_ibuf: IBUF
port map (
  O => data_b_d(27),
  I => data_b(27));
data_b_28_ibuf: IBUF
port map (
  O => data_b_d(28),
  I => data_b(28));
data_b_29_ibuf: IBUF
port map (
  O => data_b_d(29),
  I => data_b(29));
data_b_30_ibuf: IBUF
port map (
  O => data_b_d(30),
  I => data_b(30));
data_b_31_ibuf: IBUF
port map (
  O => data_b_d(31),
  I => data_b(31));
result_0_obuf: OBUF
port map (
  O => result(0),
  I => result_d(0));
result_1_obuf: OBUF
port map (
  O => result(1),
  I => result_d(1));
result_2_obuf: OBUF
port map (
  O => result(2),
  I => result_d(2));
result_3_obuf: OBUF
port map (
  O => result(3),
  I => result_d(3));
result_4_obuf: OBUF
port map (
  O => result(4),
  I => result_d(4));
result_5_obuf: OBUF
port map (
  O => result(5),
  I => result_d(5));
result_6_obuf: OBUF
port map (
  O => result(6),
  I => result_d(6));
result_7_obuf: OBUF
port map (
  O => result(7),
  I => result_d(7));
result_8_obuf: OBUF
port map (
  O => result(8),
  I => result_d(8));
result_9_obuf: OBUF
port map (
  O => result(9),
  I => result_d(9));
result_10_obuf: OBUF
port map (
  O => result(10),
  I => result_d(10));
result_11_obuf: OBUF
port map (
  O => result(11),
  I => result_d(11));
result_12_obuf: OBUF
port map (
  O => result(12),
  I => result_d(12));
result_13_obuf: OBUF
port map (
  O => result(13),
  I => result_d(13));
result_14_obuf: OBUF
port map (
  O => result(14),
  I => result_d(14));
result_15_obuf: OBUF
port map (
  O => result(15),
  I => result_d(15));
result_16_obuf: OBUF
port map (
  O => result(16),
  I => result_d(16));
result_17_obuf: OBUF
port map (
  O => result(17),
  I => result_d(17));
result_18_obuf: OBUF
port map (
  O => result(18),
  I => result_d(18));
result_19_obuf: OBUF
port map (
  O => result(19),
  I => result_d(19));
result_20_obuf: OBUF
port map (
  O => result(20),
  I => result_d(20));
result_21_obuf: OBUF
port map (
  O => result(21),
  I => result_d(21));
result_22_obuf: OBUF
port map (
  O => result(22),
  I => result_d(22));
result_23_obuf: OBUF
port map (
  O => result(23),
  I => result_d(23));
result_24_obuf: OBUF
port map (
  O => result(24),
  I => result_d(24));
result_25_obuf: OBUF
port map (
  O => result(25),
  I => result_d(25));
result_26_obuf: OBUF
port map (
  O => result(26),
  I => result_d(26));
result_27_obuf: OBUF
port map (
  O => result(27),
  I => result_d(27));
result_28_obuf: OBUF
port map (
  O => result(28),
  I => result_d(28));
result_29_obuf: OBUF
port map (
  O => result(29),
  I => result_d(29));
result_30_obuf: OBUF
port map (
  O => result(30),
  I => result_d(30));
result_31_obuf: OBUF
port map (
  O => result(31),
  I => result_d(31));
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_36: GSR
port map (
  GSRI => VCC_0);
FP_Add_Sub_inst: \(FP_Add_Sub)/(FP_Add_Sub_Top)\
port map(
  clk_d => clk_d,
  VCC_0 => VCC_0,
  GND_0 => GND_0,
  op_d => op_d,
  rstn_d => rstn_d,
  data_a_d(31 downto 0) => data_a_d(31 downto 0),
  data_b_d(31 downto 0) => data_b_d(31 downto 0),
  result_d(31 downto 0) => result_d(31 downto 0));
end beh;
