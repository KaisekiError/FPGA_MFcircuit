--
--Written by GowinSynthesis
--Tool Version "V1.9.12 (64-bit)"
--Sat Nov  1 19:50:00 2025

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.12_x64/IDE/ipcore/FPMULT/data/FP_Mult.v"
--file1 "\C:/Gowin/Gowin_V1.9.12_x64/IDE/ipcore/FPMULT/data/FP_Mult_wrap.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
m2OFuOz+NHJOwpa1mMC1hlO/PcHHENhEIqfLSbUYchGreBgaJ7gycV2D3rTrj6vV/ya0uXPek25d
rVe5/5TUTAhtEjzfB3CDliK5x+2zbwYQ/aQ+OU1Or9U7HJ/ZMRpqsamLAnwfkrpfm0osy+9xnpjP
ll8EI3Epc6w7fyw3VFTqXZ4NHZ9UrgBaM8MCyiTSUzccI4olsiNeOYFhPVxRL+A8xR4Zo734qEjB
LZKn/egMW563iqK7+lzELDhuNrm1KS1WjFF+vK+BZTL7A3PuQ0DBUnBlsnA6ua3pGPJ8fGgmJD11
3VThCfkVfRyLy3ybvp6LRASkhKNV6zLyvRUYaw==

`protect encoding=(enctype="base64", line_length=76, bytes=163616)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
kdur4D5dyd6DFE+HGehbFM1BmZLEjWc95FuHgif2gCrYjz23w1Cr1d+ZX8GPmBGvzLysjGOrun42
dUYSySmg+RGC7DeD85rOq5zEn7sQ2ZqfPDHxivDIddz7ndHDiYcFk/eo/LtCQkSQ1wgP+cVIBZog
U8BiTbVTVRGzkYxDbIdHeGnkx0tLGOW4Qq7BqpgAqgP7n4wBbcXLaj9ieNrtXv+YDaUXWCnJOXOz
R7vsTygWR7kmYQ/GNATpjWTSYyY1LtKNkIb8HN+RFZ8h8C2q9DpjOD7Vdfg8AVgye1wHNoKlDR2E
2YbE8TmSbdYVvj/H7E2NrMWXDPZpWkJOca716PpdZSLLBGKkTk1NJBEoJV4XOYZFFwOXIPgZf+k8
1yMZDKvVld+WXxZvEd+/RLqBygwZHZYyDPGxZ+RnZwI1grbaNTLSH7i9Pk4nI90TBitDJc3TQzcr
NOJvWVD74/oRLkj8ajRPuuDDPFfuuBUQ0zbT0t1u+ekDOh2BxxCnGuE6kW5Yq9XwQwlpO7/url+b
wph2+3JkoBUMfe1uliqFMOBO8DQzDp3+gD/rkB/gQx4A9mbsHeIoqd29LdUP4WX3rnVebTL7mvDK
XFk1/IXnJiRu7rn0t1o1Y83AyzMREhaTh7XD3LdQ1Zi3SXA1UKwsKWt8foC9wEC3QvXKUvGt5LYk
sgOjUQxY/ZvLMwyIDHQCxSrVS5QomcHJBHW/4veWMMh2m30MuHchDXFYbZN9FzWd+b2Na7U4BgxL
vQo//PdKZxxolqItMMVp5rXh6GoXiwY1t0hoiU/QUCjm9cO7nkKCc+3GtlXbq6OdPdMHegvlNZ9B
SHww/qsnxGIAbHFJL88M9bnpl+FtG/mSZm8AyjNek4goYJ+V7qp8d81V/awIqbwgaj60o7KAh8GB
dbExxXOgZL4TAGlHsCbdJn26fG0gJwOi8KazF/GU0CLXTjy6iXvfu2rjfzyOHt3mhRrFh04SM4wG
QWxAPtnTtY36CfCbh/zaIO+PqqTJmEDwjWMBcE3fB4QvCqkxL24dKUCME3eVH9zUFX3RG6pQVmU2
NMKElGyDULSamHLhdCUocBkfz1pBoJ7X7pYXBF2brWxiKuxrpApzlH+Y/gelT6fAm5OqsFwTF/3s
0vPCDvCkORiyxfEQaI8aK0CSLNlwk8i25avXVlepFwHyUIDVHFXx9gtM4+D20BamCgXQkjBugKhp
ZW3223dgWPJPSWtYizgOlq/5z2a5eP5Qs4r3QRSbchD+sFHJBkdx2Ezr4msX9aVQBpvA73GIakJH
aXRLnX9TTP0v+h/JXLYhCaGKgy0MUFvo32fJa0icXT33sXUgoZ0bjeLdJCuif/DPd2mHwx2gWvBX
/PhYbS59azhGPt6jiSslrC9F0Ly2ZFDF57nG74m5z1lMAFV5XPJI+toR0hlSaIZfedItfgpK2Ibl
+Z0LQpj+WRzHVKzeCF7qOMwcWOmIGWkpjpNBtD8KkWTlZ4U5IfV65nrdpmQQwWMw/f3DNhq7EcAT
mSz82LNeVGG78cjKwlVcm3uDu9mNggEexRKsN6cPORRKMgSSba+b1jxApGThw9dWq5tR8etwct+H
WzeXfSClNwsV+mn/eiDCxVh6UiBYsSfjmAmKyehxkjP3P5mmaS+yfHN5/2mtY0WRbEZYxF/FaiFi
ucD8WSYoqVO+GWHOiPWh/ApW8hZRT9ZBb/h8yVzQ/3ue01GDS8UO6ORL00xw4XEaOyA44oB1XMpy
pwnojJUHQtwCgaLrK/SAwc0kT5HbLxFMLjg8ZE0WBKoyr7eqjd4LlmKZDgwAyx6Cy7Mjy68azfxY
Sc9D2iEe4GOCh+uJ51VJN/5niaF6PITOIJAl1C47uOmy7RxvNgNH0j1s5NMjmtUeSHzGrqUK0C3i
HJ5DTdpD+fQ3/12+wG8HkcPa2w03TlCmGezZ97gWKBO/kYWNC+BPz+U09CCtm82Cj5dnOV0CpWaY
N8NswNMq7o6eyqKaOEZZfAZYp3jl2iE/TBzGLKUiAVY+4GmlvT+k/TmOP88UaT7jMbTVSza5QaiI
s3jNWw6KzyHLSL1S1e9/fugC0oaRT5xkdNFwMMOszcHV1LAj6Pr3N2Vjn9bkTDaQ692OaoDBW2vp
to0nz0pMhL8lHw2R8gNQ8A365z+4gP/TsBmd6SVf9d9YycF/Roi3BohePx5DQONcqQA3rVajnOpb
SRo4k98nvHc8hM/gEY/PUOBP3nDq/0YI81p7p86di3QDyKsjCf0DWXILkQa2Y62gEvMsSaKQBH0w
BumFTlXqpNX4rpIWFRp65o9G8M02WgZKbhI2GelMT29SSBPjUT+Nm9yJ6vu0/zNcUK6nia29Qeug
uwlUFxG0d9cNWKUi+S0wIwwSds8YVV9SGUNy3G3aaERenzPPSQLnwKwS7MXllUnu5z/WafK/QyUl
7UkFxA2ijZXxm5oGHlnCwZpUdNtwTiFKFJ/cgQa3EM9c7XwncJCycVyIIrxQrLhyjr+MYOh2M0io
xsUL0haxAmaWkeLVAmvZ5uqPNpRd57aEchXJcO399ztUnGdQJfD6PLIv2sHiI9S2FO6muZQoEzsB
tZubhNF59kz23HK1mn+JiGrKSOcfXB5CAUa+lhe8taSFkQDrnpI9B9uYIC1LbUwT3yLXnzt/H6vu
KkOs7B3Kyezrgd/iKhplXMx9Ayd7Kf8JxNRogOkjAUI+/fvrkLTGH1gZQOdil9Q6XUGLZl8cpzK9
+RvQo2LM38EqGRLfHRR365qW/t/1EaGwXtGjIMKwzRwcW40dg0uj1pQAhKR8mvdAB76fBhdZPQyN
ho0g+HMtP9q3TtPMhDCqO5K5ffD4+GvfmbouVf2OaIMGPHrABr3e3mqdUs4mmiwVy9xVQv2T71zQ
kUnBju6Is0007HUgXB3gQy4rS08B5b75KrxtthRov14h0RSJZKLe1q6fPQAl+93HUAKWhIB2J+3w
pruZn1Qms6zZraNIswViYvaPq44AJhhtkYfMDa6tx+FEfNEBhXijM4i/UQcNubCyDOBCgJp+//aB
RGwe2j5Zu4fzT/2NRxBeYR7BnWCwgXHFy7G3HNg84MnOPFlAkqTQQt6Sj9g9axEN56QlLMjGL30X
62GChcF8kiA9X3y5rDlvgZkb0yZseDKcLH1ulN7rEQzj/NXBnqUZ6/cQa+9xjBbRxqYkbu9lXyjM
KjOA3Jr3htzdM7Kq3soINLchGE/mJPSsriIFwgDFtZmQNvyCMzflD4ljCWtAqY+B4VtdG7LCTMiW
0p10R7Wl/bw/htdkmmvm0wtsvK8XA9/pocKc+v0s+WhG3wLrr8iVU2Jf/A4o21fP99xb0LgoGZ9i
Qm/weibI/lKnAhtx31JikGjaPzq1H95WnxssTysPrDdud3w9RZ+kHdF6cqEQVk/iCLAb80a6VHKM
uLsjxQFb2TkP9O6J7nGFUAhJaL61wsYKCzOK63NNmK0WXfeoR2M6l9luGuf4q3mSatGbfcU4J8Og
B2MgIRFh42d38vGm8YzIsDRn5SO+VsGt7kEn81JoBqJRiuA4dPm7ZKeMV9nG8Bzb4rN+2SE9j/6E
uJca9dxFXl6pzradTyyiaV/b0v3wy45xLj2rYZtnrILrBkt3GsoqGk/Pm0L384BStpOPOX4+Sj7L
IQXAfuVtM33eADZ4fd09COOVYuH6dcrecnAib8wMAbJf8mh4/8GKicbTNJ/q3s7XlGCx65kNp72H
/kfrYDWDI5WKVZ8E6iStNCsKhj6qoD1Xys9lNo2pDps8uJyDYFHfuCcTIFb/KIP7Y1WUfihRplEk
rc0BuwGCzowkr+iDwx6rm49JuQsqnzMF2YXbPz+Ya6inBY7HkSmALSPchl9ILKldg/IP161yiSpU
gs61TiUSbYuFppz6knvt+k6RvyxcGbr6Rfhew4jsmnRacVJb7bwD4pfwAfe6ouF2/YqZY7SHsV10
Dwe6Qu8nUe3CPwBoSx6AQ8dEgm/tnx5k7ZazxwW7Qc2c5uPX8ZMfd6wu2fAz621gAnQGxW3jYruO
34XhlEioVxRPhuS2+VfQRLrR4OeRevsWPnXh98tuUOB8b5loNd/7v03EQgJy4cNNZgDV2ACYsANl
iH4NxwzgLU48ANwjsWq+3x1971IZsefOwHfufZBRFHKcYS16krd5r8qTOrCAzUhqWSEZU+r8ABl8
DGh+wwOTVun4S9ZljseF+2cLTM6oSG1qudgIM21n0EaDA0xAFXKZWNioUavDmFbtb1SHCmzVAqan
8vjAvrzw43qRLwNW639alNOUDVxN6C041c26GgJIrpHHGDf1lAAySNq1Wybw/35uuJg/t0dIlSWJ
VSHk2liZbysPBkRVSlB8V8mHGUd5UrvcyZ++UVqf2UDFhSvgHIV8lea2VVNEtC9+R5RLPFtFrVar
cNmld5pHtH9whr6WNeQp/K5/15HaTJskNKuLz7MjCQdy4L+IkSqCNnKOtrmPp8/ME/CVuZbTPnAn
CKBXMpjj0Ct9qhRyZ++rLU3AfPjv7eYw9eKBNBdx7CyjYuio5lbZ96DYjNZaksxQVn9nsuGFWkhc
Xi4YxmZqqtZnHOTZjbYdv7cJrSDXvC8ytntTN8x2mAZE5O8ElrysmENFHzeJWoQsqjvEaYoaDqmr
3lCe44FDSIwenld+uP7Qn4GlMjA/UWiVZUsE5sZFhFxPk8G5LTktS3HDvj37F9al8ytoQR0l6mDg
FnnijsyYvHnuwNA2lO6AeIbxU0j+ng6cGq2WjDM//zWzNqe+pi1Gwv+PWbfg0B8WP8o7IDqccPER
+Y8mcgWaq/H/sdgGnidGBdTlB6tWsER6RbN+RI9dr7uHe674hbUTsfECThOxxkGA5/sb6l5Me+nB
izk33G5LCnd9fQeJBRw3r7lYmPC7LRZayNENNgqD0T/MIHJO1d9mBHaLucfbDQ1O6JTzSXr1pYtX
fS/AsJ792sdcKkQ7x0ds78nv+hZ418FtTLw9EmtBoVgH6KK2RktnUd7bplAoAqFa3rG365WTKZFP
Jd9ZD7qWHEIyMo7h+JytrnPJV0wvkWZvD9z7YfcbIrXrDkLfTsxDS4u7Cw4OB6lUQhSeyHVE8JJ+
rC8Be2YoKOp93eG81OOwQPjk07T4Hqwc0W3VZZmygxnfQFrrUOT2onnxeSuwy4bZ5DvkQAjxchkF
dXn9UOY3HN4oMMzi7cd9hOgFUVhWiTUXNfxThWUyXyCNwKgsCg9CWRMeAAicEReQZE8Px2X7X6dQ
C8CflPSiGuhoMwRueThRrCDwRHxUbVSaG4wVp13sjBx+WJuA61fclUekRoihu0TWHEmdUBeO9tIl
M4L0XYKdudEKxazpQVGN1K3lftWJUmb4XbfruS8LjX4Zw+TJmpLZQAFtIk4uPmHz9iqiaCcRuMhe
x1Js6OV6ldUvve9FTrQ5XVfiYhG1mieQkStJY/qrHFPTD1acKExaDmSg083CrBlmNn3N6r/jYn8U
L3w2JlNBR4nYrY7MsyDbZHec66buctavXM0BJnLG22ivMn+30CVrXTkJpLDYzEoH0MmmbUiINFk5
EJYpEzYM2OkvHKDBv2rCeeMCeWSWoP71iIPLQ9bU4/BeS2nVjazBeQCca+MzqAcQkwMnpZwAIzpr
20IXgnUB3SCzDEoEpJQRqfHUWdJN/U7IaXckRNMcJEuxAI9QLERDhNMy5yZHOrBT50mgo0U8DR0w
HoYZBaunKpgZB9Qvjl2ncEIsqPuJ2vBxqnyN2W0uzFx1yLSoRHpFX8PMaAm0dxO1a73X1l65N1Ya
fEzG5MzK4ipsJHFHbrEWzPyDCU01MYoL5gNvm+Sw1jrU1uxRRzSeQmcdTjVq86fBZ26e+uVU7qa7
h+dsdkXUUW3HSWb6z6O1DMlmpHKiCfwov4LW0W/mbEyAjwZDZ5NQStH9h78sKagNzp71JjUHYryV
qLcfRZDhWAMH4iO+HfzLcDo0ppPhTyZNurmhUPUEDWF7jTdTVXq7P/Q9PXPF98HCIslklYqkxdfh
aRa6tnuPX1o7hhnOhO+nOFsJeTJIvT7jZ/XclaZOPE/GwmmEd8jGRPWKi9LKv56PVDy0DJhQGXO4
4af0hnLqQFiNiTsROCGJ5CZjdQz4bhVFxs4BnVc5GtR6z9Jv5GF8gIRM/hkGkbCN+3maVJFZJ6sL
DwDa2DMdoCS/JSuRI9zLi1z5wpw+WcAVWYYMqplL8gHMpy75DaWg7pO4xxNNIqaxY+nPRKFqYy6g
QfDmYEoPWm4PKUW+wZGN0O2kQBoTtmAYOIl8bJDFaTk46pJb+Ya9T6CQZBdq6+7ARenGz3JHrY5q
g978Dpkxlql+LNhiH6eFe0mP8iY+nPlTiTZ9tw5xNcpSMJ6E0rlhZ4UgpaKRUUJlPuBUgfgs7O6u
Ox/O9fh1loI8oPGBplobgc9tBRjLjzxmfVfvmuJKE4q17bzEBMDhADPzkiLpaRHpJlT6I7Wv4lGR
ZBwQwoCOVEy4INqT46RbIf7+ln06eY1TBEdP4esQBC8E1B9JenfJjwMz9zmEcmNtqGozFygoTMvI
kZnFqUH73iV0fCSCT+AyiBKyG3N0qVb3XkmukI4l8fDFxZOTn65C41c0XdSgGTG3lU5Hsgki79Ap
ixgYQ4K1ZacGX5cRMTU/R4JPZjbly2L1wQrHhcc4gWTqgn1qp1oXdQAxE3bOopZmcdroJa4OEQmV
at1AiL0KTbQwEZ3Dgw3BNRTtC7QSAmJbPn0/SIPeK4owBShccqO54S+zQk2sjWfJOdtKS6TUU/qE
RD3HJ04DvsLgA0PN0mb9mOCJxxTJMS4nFMqC5Bbh7g4gwqvbjT4i02T2W5LmMqyAbQjBDz7sDXZX
1qpNw0HC7s20UaAlM+zPKYoEvO97HpTS99TvJgBOEaXAIClzSBgzqegDtmW/HKlhtADMdsIVnjn3
PUeO7s6+3msHAO0RhtqpixG246AM9wDcFHEKmXd7XQIl2tM4ZCAq+jOWFa4/tFGAKZx2i2bqFSvC
zFPsg/oGf51dqhTJZ4ZYfXdBH7hgYoU6fcf8ffu+YMbHVMSt0I53yapVych92aakVibDPQkUH6hV
keSmH4HN/Cq4hOsTlkJOS1Ks6Fqe26oi3GslPDrJjgQrajDWuPl8KGlxjC1PXasIimxTzjqOFI1G
g8edIoqNdm0/b9FvMXIWhFIUZzqCoyKVlz0TtFm4ZpCVH/iwXGIjQRopGbc9bVbi6kDOPhmUpDGg
q+Jw1GjgAln+m1VaAwdKk1KnDnO+gMBlumpXjLJLadBE642kF7MNAFKfCoPMTZpqpwofYA2wY/HD
t/c+1lNs3k7QX2lXu7arxP91MY26Y+3O4PGb4el8vab0SnlWP+dZDVTLO1+ldsT+5WnL9l2w9TUn
NS8fNtJStqngiGqyDpAU/iemByPxAZPh88hL8U7zn8mEwmeB8IVQ7W6BDQHDcwVOSYfnIBX0H9T2
Pa+Upwo0v1ULJEa98/WgFFWwSipEECqSBbZ4M7wVcokPyozLnOMw4U0Kr6rHAedXlwo1m9nEbHD4
yaaGnstIdPiwrS1C6prAHPCbvk7jY8b7tpBzwTRjKbMC41aVORoTBt3Hw/uupWSKy+macjrFc7g9
dwjeTW5/bPJNTcedlCzLJoDXVh7K2r25MPkqm5fnt+Chen/OEzig3z8qOD4Spw1NJPXgnu1wTwUl
FIXHcrHON34gJjBqBJiwxy5W3Fe8GzJ2SIUkqlTSZ4rKfY20mgbtTXYvFawFERgGl2tx0IWCIPQa
mupMtkNI325szZZDe7nDRqwJVobRtW41d4OY+qfdKuCEJv+PH1S83ZZ/dkCa/Q/OiALp5v86tXU8
iYsuiWEke4lERQzHbqJDktV8kSqaLIhpLOmG/hQkgfvUcPDsSB4J100LjENXQYc3uQYEcX8/xfqA
KfG3Zb604xd4NsMxivF3YfaJLjJMWazx0uzaDdz4GEV+nU4d7cxR+5a/+6O18i+nrm2e0jH449rM
nLeb+ZU5hVkGkb48/UXRHdxzgom5+Jr2lwxvlCiHRC2TKM+U9q9C5IxyUejX4Gv6a+wTiXnr+WoS
xaR5ZswKCfWGcwGBk/gOBswFjg+HBWT3QYm2Gfglb4xeQvONypKunm3BiGf2INRj7S5y7e02i/YH
Dh6FHfB9Lz2eaqx99gyUyWf380WeNxAZPQWT1y+Rd9QozaNLMicgF7OedUrFncqxA70AtmD/Z9qh
kiHo+TyqqfEcnpNn6Jd1RhX5r+XxujZodXYBeVsWdWu3FQi3FNvz8JOP8elVOk1G7Fe4oRL6DG/s
rK+0XVydyTwMEWUOyoDKXzvnkyZ0Eh4U5w+NxEM0CXUuIgH6UbpJg35g0uNlWAujC2SYkPRS+lcP
4FfirpuZ4D0teP0JmGd52P3LtTT4xQlsKSk7mC8whC8PDIygGW2N74q+MhrZdYcJeJNsPdbkE+3y
W40ClbzC3AFw+nCOQ9zCdtmxJkEhPTlCt24T3uWGw24ol25+WazzFPnyOgewgDrlUWMn1JljEaUO
K221LwP6G5reK49Gg59c527QgH2pOMvN+41vCfBs+Gv7FpZUvoBL1AfpaVwV4nYOxlHpp99+9AgH
CVdZElOAJa3kIrK0pOv5wipTdCMwlpVt8Gyi6s8tg6c2JS69EqHSe0xARLGZ+0rGCLGWIiux2uUD
T1E4HdVAIG3myBzVk9Gv7FgLlbV5n9dw/se5BpUu2Ns4/YqUODJ6/3Vm+zgOmZnEsKAWuVnV5maT
n5UzJnCN/YAZWqEz7uvQ/l6nbjrG3w8i7aoM749wps9OmY8yuxMGe0cO0BCrfxvpcVAkYrHKI1oe
Tc4dlMFoGalFSC996u0OLkEfumgk6NtCqjpqK7HCDhrv6cKTzu6ouyJeDcwZRaDKQB0AaRzriQRD
KZ5aDBRTNl6qGVEVID3W2AylX0qO6uLo4TjJfje3XdeArVLHOfqp9w1z1dR/Hr+b5bEkLfR12GYb
LP6flhmWznrkUE4+9YS1j3YfpySup88dmF6rMltlo4F36SLqg6x9UMTPGTdB2gJJ2B3bzfdSs8JL
7+1p1ivvsMXdl9xP3HE4z9rwgLDQKWohR1K9GWQ/zI2wI0YF29fFz+ux84qbE9GI7re5OSrD63to
2zkS3t0NtCsjxEF2IBMcbMCarJauIbfN0VotwIAYmMNc2aZBxC6+O7pYjG1dHdldcBYCgKKBNnW3
k0DYSshaFzq7QsrGzaSqnoMiofHCXbYRRXhriz0HvvmmATKFWyy/6eqXkqRfJoGEl74zNmjnIrTP
qyne7Uavrc3sN+1Gnuq7M0QUxmkWVku+P6IRWsdFbt37rPUstRJ4tKMXAyAchJWipdCfD1x3bbhs
SUXDp3Z3Pj9vJD3N62lcm7VSb7oEjAn7Q1+HgaA+hQL0SNFttWvTG8qAT2rHpWHMDJ+l6/NmQzld
zQ5cC92+or/PAdTqq1KXyqJo9fSPN14iEFbWdxBZ8HQl7Jg/Z4fVKSFzMlTV9ExV64cB28gBDxKY
8sGK4Qt1fMc5zgYm/aWkA7cBmzx5meUZEbx9IxujHN2bvHppWrXSGNJcNvVMkhid4ntroB/h0KyQ
PmCDeDosa6MAYg8sCXy0cuIi5DMhxtThYd2TD2JMRwLgD8RkUFXH3ESOowa3JxFOLOY8MEpFOLcF
UwNw24EeLR/eqgdY3CIhi6xRb+SYwOjze9+mzXpphl+PQAFbbzi25CkH3PMf8nNG6Pno2gh0osaj
75xzKM2BWs+w+sKA/2S7BYwNCqNfwj0wtpxEOjOW1wEwJD91E/aJQ8g52QtdasaYFJZImDB76M6T
EnfVV05SHWTWNmZOW6JfBJVrPj6ujtlD/42minPmR3Kdy5/qmjhw57Ptj143Ofo18nGhKOVTu1Ay
y8tWgDuRlAAhWRBKgsyQVM1Wh6oNoK9MQRL7tr1PaZXaF7puVxCggqF4U2ZoA18dAxIFnjQefIFs
S1yvXyyWId4kH8YgoiBEif5WJbqrtDHW8MYShLM1rz5PyY5T5bKD4tTQ2zfMPuDRhRuVbolD5Omz
7ddHLgsNhUCreb+51xdEC3Jl3FCTyX/h7H4wubqBV8ywtOnODhMWuA/uDexkBq4ujEAoUHPU15uP
Ai5glkbBVqdsy6okRqlo2niFcovvvQ85PEIO1z05VajaeV5NDhsXbbr77P3Wn96rnuM3HiNglLab
4E1hknAe4FJu9jP8NsPPVUQz/qlrR4mrpPcLIluGAAQbpfiJgyZo/p1jyk3DPGF34HYZJqCSoidm
7u7PshiYNwMu3B6aI0quEtTYmkeNy/hEMGLTtGOzKs+iSm3RPIo1xAFTa1Ew9X16Wx4ADwXjQbwQ
cnUCMtp1W4WiLh/52hpWKpiPAu9OPOgCe8yPXOpdL/JhMDC1u3rGSfwJGmJ2pekSi5dnKnv3ZHV0
49UOKFX2y/45E7opdLBMtG+Hlh7FfQ7QiXEWuVcBVpVEHKvKDm3/Z/mL3h2OABOksa2WM9qDDsbm
LDJ3KPNfkzi7VblWKI2+OuwI4unG+tG5VG9DrSEdB7TFzb4ACTFD2++9AmyPWzZwOL/g4b43emWV
of/Fq7DaYRvBOSfDx5g5Pk5B1hta3gSy4WtjA/KAXsM2eeDOuFfpXmYjChVja99uz2Y5KDH2cve5
YR+g+i/+6k7NmPHo9Ql3Iz2tBTGpJBkq9WkLP3AgCPPf3R7v/mvqLMiHi8sDmAjsr8J/TWa08Wn2
W47KSuOh1Bqbko6Nc9DrL2x4jbMlJdXScB4XeebHMKUXIudddFnQvM3l9SXCeuocImQETQIQjd0T
hc2gzIPoQbne3dktY1B/4ds1Px+t1K5iSMDxuIuSPf4rl8fhk8Zj6mLbfhKSk4sBuYOHvqcieh20
0A/X9MdNiR2fgRNwWGsOt9DvKn1QT4H8LSG/175rD9T2IEWncqvE81DMQ59Uza9EKR7m6k/bn9jK
Z5bS7OGCnDNq/4h/NoRYYLfIceIchVyY9tuG+8nJDhb4h1bljy/nxrGxt9zGbvxKTehE2vztmsnr
hE9E7p2ZAfEAIfkGH7iMKZm/vH+kkMeklEJJ6j3meE+rZsJ5DDM2dNIImoNogeL+Eq5HxXWDGF0C
iaKrkUuKcC3LuHjk/mO88OQGAzJyowsYMer9aAZZTknK0kXmuOpANrdTdNXZMMx/5xJ5FOVWS2X1
85yCb1B1q8SupiAmTe2tq+cQKGVG3MCPhB362TqKTMgMgFnZuqO4cOuRB6yv6sZ3qQkO770wRqU9
Tk5hKfK/INDEehzP9dua/HBzaequHgRoJQuJr4fMsCx+DroDeUKR+RhI8t2Oz06L/xQwSMQZ7jVP
PiyCS0hr8US5d8XfLEbFk1XAYIRPAZHQ1lSdFnu46VbvVhoEE/t1SaDcbk6km+atd+7/ovg8drq4
1V0LfZeeY3siaG/gSnfS3sTjffY7ynYQeeTcc8I4MBcHP36VFsvykm53Er22nJrbmGEX+d5+VIMQ
WIImXKhOypOOoQvd3KPcqycXNDtPmPlY59MkvfURkYXgZYESIcPpDddDPCvlCNR0ZiSgJna1j+Y6
28pvN/8m7CyLW7ePzZrp53gZNiDcSxdQkntx4+TffuxWr3kae/Kv0KmLHAKze3tg8bnDeC8rksUH
Ux8XPnvy7lzjw/q0Ye9+EvDKdmDF64YLjvIzW5kGGoJ3As4OSGB9Ux1YqX+8MBqAGFNkhSlouArv
Wj1C05SwCYGEDbX+lWuTOg6iRHbP/rI1V5avXogU1++MRb44v3vbao+UY0w5LYqrmZTjFnKbut5u
4EYSf3C3zbTLbHUTnKx7M6jUlsuPEQzr/Sqz0VvHgPOYLDfnY1RlZazWWsaJEy4vG2VwwEhavLEN
9q0yy7iww+2EjgPqYsKl0Nziaou99brKZjMlKxhYgQsDeEQDHZDJyF7R2ypGTlMPKVmEYordtg3i
R6FKvqb0s+7BN6O+l8GpO+gx7cnHKOthSJrnGGalHLtw+y0vsPuG6EwzTMbEb40vt2JxuJp+zxyA
7QTXQZCTOSyMxqhsQUNkyTHecjlfh53MKfwt/oQJROLZIaEiXt34Dr7z5Xt0muwKRCzaIIV4iYqC
ftYxj8P8fsNyTQpmVQ0q4u4USYYJVbHItG8RBB/ZITcjOMpNNGF+kqjrycFRGOZRWCtsGUem1M/O
kpw+0EoPQyaOe4dzjPEtAe9jPkEyIZIiEbQcsi9qSuMe8av0d5oUqD8hwjG3D45J5CluTWwSG2HT
QmDEoTZsvXnavNifUwJLdDJkoLre+Tl30cVtmJ+F655pFKVrY6Tmk/WuJvob9yqY7G7+6mPGqdQv
U11cNWI/D7rC2vPaSY7z/TsXuKh9ojT2fT9p6JqRFOW1OdsvIuGlLJOZtEDh8757YONEIKn7PYIg
0OLiM0oOl1avVnUsrO0ZSHYhBO2g7U6mqUQNcgsJnQpRBT2/qr3gjviRlAYgaS0C9NHPnjJWQqpZ
lM1gusv8FFtRpI1Ht3LJlTfaQP0IVEJ31V3XCSqd77PUht5O5ktk4KywEmytE+bzSvXsYD2LkHO3
gIEtslgmJLTJNp6blToD1nY5aqIZ2Sl0/Ud4nP471dq8kRtjNwlXwRW7rn/ovq7cu9y+bxgL8mLR
ixa/9nloWRI7ue9+Pl5Tp9gyFN3H/zpkHJ0I3cYIEd8GnlYgptN62RYCt95Fq+BRPtWenPUPqp6w
/S/xcLl/Yrea/6wAkNVHqc4IEONJ34ILboAtPJOGXZPiN+HVc3ICdyVzXEpHg8TD6UYOjZA+MzW2
wAkG0TG5UauLyK9GNPYbXg4EJJZEcPHyJCSnupUPErNKmHWkbkkBLr973M0xHeGIvFIUdn1MKKTo
hghF3eVDkYnKLnKMp4eVEcnZ2GcOFpoVuRqIorWwelh2rZjT85iwpH6Y4U3SIGpbObvIaMgWOfFv
If7KE1ERfRLSxSk4VbS9SQv6ySzi3ZDGbf+GU6ZcsKb/u18sGE/LVajnpzLqArPBPsrLTrR++PGH
faGj0BlLcUV6JNrmshY5wtaxsigvYC6bMXxq0X1EGy5ghFCyPcAtrPx+NWP8H86vaGy2U14mxKfQ
cWfGnuuiBYW5StFsQAOqmqrFt88tqIcVvvGfyGgSbMt/xHEr+wotqJOadyYoLwu8CWdLyS2X8mwe
75GTSnjzmec6jisHI66Z4vxEL+1mmjkoxkCXifq1OXHCwPDzKygny1eEj0c+Kc9DvKDs+H4swTgh
Q+E7l1FATaXLfiQbuCg657LX20GGqOo2oDGBZwVIjMv55Obqb09K1RkoRPaqt3YlJZw94RQcXB/t
Q3KpeXZjnlspv+Sh4kx7rWhZDfNvvVwTZvfAB8x906NSKOT3p6SLIBEsDs6lpU9RjLbOoy3g/9B0
1WsSw67EK7bWy2MVQ937jpDT23kYXrw4vNlSAuQAGLVpkOoMopUN0fmNdOpyNAa9kPuP5SlWsqeM
eB4dDdqygx4YVBWoAwTAXwsLfkjq6Hmw+Bw7FisX73Co2Xq0xciaVgVZgYHZn87AvBnlQnChJD4o
DNZX2+/rvGx0Tx5T3Gopycpt7IdMcsH0DY5Lyg3qb79TBTWI4+ten5n68tplIWj9Zs7Ksf2/E5f1
k/waqjWDcf07HYBxBAAOzIR19YC8e5mksTGQ/U6pUU2ERzBXLvUUKg+DahKiURYeNK3U4UcJSkIj
eHR7loIPx2LUIFXKIzn0Jy9Kemo9XAjempP5uDybqb5LW7SRAWs19lNUJxJLfUcIXmquX+rE96a3
Qsk1vynM5NjYsGsqOAzYoF5gjPL8fDGh7EwekURSIHv95J8LVDMmNVMQP2vIs5z50qcJfBdbunXP
pIbLq8WrciZZJOa6p2GuzAcrSi27wvQ8SbAzCG0xNfAqbRh0ye5H4UrF0MfFqg5cITbseqVLSltJ
IMP/12WwmfdcKI+0va496VW/xP5tKzFnMp4MS7SzUKpimVCeD23GeQ0wOw/BngRWZR93wxOnQGv5
/jAagLj/0CmIQkMT0/d7ffiDAU8Ha5rTr8CwxLn18PGBFX/0EkDqe5hUnNX1tHLpifT+jaUJCcIL
6NeUpiE83+BcnhjssGz3d1Vy39n1Z5a0hL2s2IRJRBMvTK3HXID3JhzgsRWulAhf+4D9PfnS1G/1
mH/uwIIPuWG498qjy/NkTt9FpQL2eu/42cbkfFDUJl9ZjRPyW41fK1vMA8K2AJ+tXJaWu17WARqI
ot9cb/0iy9iZUwUTI0KI10q7yxVTnk8CyqnVpcnyasvtzb/bSNJaOBLS9NDdL0tqqBF/9BG82Bcd
0MgUrdAUFHvveIhVEIxzOh13LhY/zLOMmqJmKwl3TzeNGnyK6scOIqw7O+udjvHSQdsFn5VHZv4x
eMtqWRu4eSmT2XFjNZmwpOKqMCnGAaf2yJqVa4ARZdh/+gTAbKVZ+9yKgOb6eUuyz2q3viwioJ31
Erslivzq//DsduEqItGYxDC2gIqPF4ylB634SVcSi9A0ZqzkeEbs2fHTaXg1Vj+VudjJnRdQTBQY
HlY4+wNOwWSmI60dgrV3g2goB8TLEPSsgwdKPxLlcT1hxj1z3A4IT5d5Eh8w0ygEQV7pO6l2J88k
iC4/2dd9Df3wiHBiqcfRMjOIw9dRMLCS3n0C0C7Igy69cWBohy26TPbm4kFMd3ne2uQDDd5j7WPD
iT+zGnEOmM6YW6nyZzyUJYDVRKfv87TswbPJfBBtf3IRWVFrWOSP+Ku1JGxI38Uro2bC/FM1OUKq
fsxfl1UFgCFbRw9PoxZSW05Xrws/mCqVSzi/IZt8zbCWYtI3RWNXoYeCJ1S7ouP7IES6/E86wI6W
u5sLrEYWCPm3RvFO/soQuc1+BrF9mXBZ4X7h/SAMb9oivnUtfPWwhr5NsxI7BnYL2tmA5eY1hnhA
HVxCy6NeFXlkU/HiE58a/BB+ENEKSeqm5ukixFAFXxVhkwEfe58StnnK+UIHePG6ID0Oxnimg0Fd
+3vq7AzS6JmxgsUoj/try0ihcnLh+nOdQ3z7i3nGyZhXOUTCaZlnUCbNbZJilDyMSzAaAygVLWW4
KvP2XWpdrLUetlGymu1DFCKgxlcaJmTsK6OHmvYz0nnppfvYUdpyZxScEDmgaT6LrxaNHrJGLjjz
HJKLKRx5sLzg6hvspjQdAUib7XGfCAHu9TaXEcuXy/kfYc3s4DO5XlG85grW5z5ETq62phfpnnaW
3u1XbPXteh//sOGtuF1nawwuXMbMSP0ozEhCp4IuRP2bt6CCqljvtcdWZBk/9KwSXDPuy/biA0uy
rztNE7k2dd2645lrVNK2jU58L8sgAi577/UdLOBR8m1CqMu++5f0907sbB2AJC8tBB1yl2RTtiIz
j3dzQEGqldUd9gYl+WYjWxHhkJrbnLIUyfbl1SdKDtdGcok1x5adrScX5AFaMGqR+hGgvKi/8kCz
o8wHPW1N6es6UpovBxvn+AkPdt9z/0T1ivVmNKwPMaapCApEQr/DEjkoXshrlSWNGw+7ZG+J6fUi
oF4u9SvxRo68GQtoC5/11sJtulxfmByTzfoR59uv0CSx1z9ck3FumG73QfciU2A8F+n3dS2Cy0wA
jz2N0z5M8OPIVgW5lFK3o5xn7lXEDRgpH+mx6wqxYjmZxBf1l7B/zT6y4dBWtHRbs7TCEGHmx++G
3YKFvP8E+eaOGPoagaaaBYE/JzU7gUPyVWIlSGT8n3O+RbnmpKzwUJ/YlqDOkt6171uoU3MvoTm6
1zw1Yi/EUeSAuvmtJbM3sYqPYVK6uJAFn8rJ6Ps33B1svaqFFmJCHL6gumOMuIE0ek4Nh18cnJdb
YSMst11+/arjr0oackqzsbAMMWO9Wt5ZqOr/F9X7feAS+x/hPfcXNGo0yW4mYEmFVkY7p1I9vt5a
serpcWwucfsZT7//0hsKpmXYfaGqjfA69XOC8+zOxstr1c6xsQzxajwRz7tCmalbMnQe1AEw3JNz
JWH+cJybeOgEDbanIkJdJLLcJ5GL0lSRo3ckKBuZftFrZbxZxYBnAQN6M4Zj6FDQZtmynnkeIZfu
Mq4OroBr+wSInTt2VBuFnvxrZ099kaivQh184dRsYMo63UAxQ5sKTfXNFbsXZVXCtTI/8SGxtSMG
lH8NchxSCFFszZljhfoZ5pM/Z/+DgEj/9ZhK0PVbf7GpNnNXZAQPL1gQ1oyKg86k9V8kR9gqTNVm
y6L1H10nS+L4ti4BkMyVeGyesqVii7lvT6tQmmI6IJjLXnbQssRZI5wfNw5qgb1lflLmEbuKEtRb
DuEAFTu/8kts/AZ+0rLqoKBUCdOeaog6dxDEGyasDuo0n0CuzP3symxhAE2tiKyclOj+3ZH90aD0
1EFzARVkK2LrU/jhaQ+uPFUNXdZNNDCGptHXWt9SixUlwT2YsVBOMkp8pcos7xjC8cuSVDfbwjXT
mtTxnu0FB8XiXXeDDULnOy4hlunj4m5CDNh7YfObwpZ3yuY+JADO0HpkTAw+LfghS3Zj8MEoMU/C
MN2XyTs/fJK7x7dwWuquy7hFuo8cyxJkUq7HploZA0Doamzr04a87kr/Yss+SpMnQJbl4yMo4gzf
HS4Flxb/0o8a80G7n3GpGgm6iFinfGp96pnYw6q31p329QlnGy+Lgl/BkTuBm3vP7Z1v3fxDtvZ5
580QuDu4Qu0KJQZYbmg+NSHzaaznID+xEkVXkMFeZ6ASG8zeR7rNPeIacqapTwZQr89OnYaZJKIv
lp3C3QKAs9/s2gHE8QRR3P0DCwFE0AT7cr1+wqmO8JiaMeTWaVmIv13c2lgZa0VNNiSP+Yn2xeR9
UXxo7OXCwklWXvnXnnAxAvjGsRkyDlB30zjzcvIOM6aPtBK+iCBuVpvJjuphgL/mTaSWo4VEddU2
fD0yD20977fc61xSt2M4wFqFHBCncp93KL248l1fcK0RKaEpMz9AybpBhCWpuoOv4ngjViRx8bux
4sLjo587IsWYMONX9Xa2oNK1BcoDD4K06JvXnyXbUK28iyHptGcvHjqoiz+SV8+orWw6qKr+WGIW
n3uOoyJnHkNJYbizOn0AvTh7mjGLEByiHDskbecvO0bEg6nSIZ3LoSPguu5DFE3Abvs/Wzzur8aD
Yme8w0qblRHkppbKG3rhBYcGcklafRYQXWE8ILV54X5m2y4FLIQu/iN4jVLKnx1cq84zC7ePAEU5
7MEMIBfAQaaONEC2PuUo5sp+L3fh0KJmA2+BBP6AX0E0dS5+Z7SJj4ZQG4QqZ3uL6lsGpHmZePlB
LLdnttuN/qpsOHcEW5Qz+8h0d0eaZvuZW7lIcbUNhf0xrEUaLX+LtVCAbhtCKPOQuxPs5bCUh8/Q
lrqglSZH+vU2XXSP4ohV2PKZiOBtq8b0yf7Q+rdNButlX0lTUO85OLaC0MZro9CZJnxv/11289VV
KNDoWDTkyiuONFsqRJ/vjqlD+XxIw7WM2UH0XG+V8XhYwoL7Xt5Vo+qWLPHZMY6ag2mo0GTHH59p
GYxNcEHDlw9TtdBfFUdtIp0olcrUR6Zg+/WQerh9IOSeHfUCb8o4omDRP0maCIFAB5BGqM0kmRQy
gVFivYrgwh2o3ys4w3+Iy1uWhxk//R8Mxp786yPJiEb2mMBHe3UOBrlg/MiRfpRtDPF7JtWOiCIV
2bxRBM70lkIMQGxwX6JwGy9bxqKPBzz6oSqgiAOf0vQooB52ZoJqeL5WMEr3GATptKeQjWTKwYF1
m55Luwfwa6puL6pXuX5OxWCaWTXUfcsvoOXl8JjpCazNCuvSP7rKGgukiTSfH0STNgJzuVB6YrOC
a7geK45jH547SrCAx7iXGPXXuDuyxPPqsa0o8HPx75BlwoD5kxxZmAm9/nrZ5TlyZM6oVn87yr9W
93uEk6ZUDGnz8NRKk0zhLAijvikL8Au+zaNH5VH+09cZMKUHsWt/bCLcxuVfkDHfDj9rIAco76u4
CwF6FyGJOYBLiyWrHf516r/ov1VnUQoIxR6Ohzdt1QnXBVVZjdi/DWE6FzdN8QGycx+YRFeQF3mO
SikonkMIjI9XAC9SHfImr5FER8jPEoD0APm73vMkz/GxhyjCJPPyY1V0kK6NCPGKosrtrKeBCP3k
//BzG51haMNxk0yjQGXo+o9MSMXle06qWj60B4/DSh5kxZwKEq6lyxaAyjsuwLCDANd9n5D4/NRH
kGYbZxS2JxF27pe2dPziGow1LYJvm72NblqYhf60xh933AajDHVLO/wpzpzvvIy0/W9Tclk1k76f
0hGFEm1BkJCbLgmHXsgNv7ir50+cj7/qbnjf3FHKaUG4QUEonOml0bfsknqBOZXBZ/+9Yp3LMndR
fBLYIjd9bh9kr6g7AIXMt5E2aCu9ZvbX+/xqj53i54OXppYfm4ojBla43a5jF2Q6Ue/yLPiHSl+g
2tpVolhyrO5GIdyq8kPJWto78i13Zh9TS0jdy8TxGyqjd+vCIVU6xoNHsgGcFTcO4WrYHtsg3OsM
+05xR5Ey1ASVV6g/ObSaW9cv13f/5r/YP4EyCy9E0WXr4oAGx7CBwF1FGV4PeMywFiFrtsp/+rB7
5GQe761amgW/eUEwuJn4xniwDONDKCLzw0gZMcOf29MVMS5M6XPvPTjL1MFlS64EMhuQYdN4XMun
PkJSim7RshYMcVEsinnnXqDA0j3EeirKxtoCaqOB9ORcW/+MORQdQ8Qamo+vxltuDF7+wxTAqKmY
oX2iHzRrZfN3GWja4sHuYEXhoy1oqRSTrwGiiuOOkaPuRI4pmeulAOUv2x/aw4IKHWdIACm07Zxr
mPzFXxEBKTSjT5cSt1XERWsIwCuCLDS1fmfxazku28xFfH+immLqSDuadKnGV8TPtr0BUKTW35pi
3R02yIkMUbA286k2eMaU+tNC/wug88sL4+/ETHYSqikkyiRC1DzZwnL33UKyDPbbM+/yvL8sI7Z3
TwwrtWLiIC1Fk63rVpPm8zKS5ceoRpmUj7qLSKTOt6BYVjlHMmCIHlGNE5A/HMETZsAIRbdc/rr4
E2E1mXOHf8HCT8UP7lL3rQCPI99g5EABVOS7iXU2dizSAJUBgDNm/x9rBXeHHIgOx8Sq7GS9oC5R
owkdM/1hLprJ2rB4VTvKS7CfxmEY2/B/RMvPe4wjPN1lJOvwT9+1rBwsSLLhxEMYwsg5+TbzV0AM
eOw1zmd609ch7oXp9izHHIl6zunsbCRahHFoFfKowEtNmlTVfN8aoRYsH8JZTDlo2tgn580eWpHn
LyFV31Dju4GLOW7DQ56jQO+Y1l8Y3eE9HaLnFTM+2Pa3igKsAeLDebAjJ1Pg757kpnTYbwC/VVCl
3Lzf0Fw3Y3tfAaxvBlwUzOL4ivflEMVJx2uPpkgNfDzDRIY52bXxu81YI3wkOVbIM4lTecyYoCC/
jWwktQH+POt4n0f0fbgrhXm9wsc+LtGKsCGiTfn8XOUJDDOvadqp1Enqn8mQC7237WN4XiKVuVBw
/HKLTDNySh/+g68s9Aa4NkFamo1xHrt1Cf7V4cwZpg5ngTlUz91idm5OpGHRbMcLnGP9vTWY28Yq
sPfWD1jEx325Fo3Obc3C8rvwc459J2mvbA7OaMOBUgZ9NlE+0npsfED7Q7L1A/g5+zMY+64fAnOr
FlY66uVGeMubYRhXqKq62Mye6t2mK7W4zC+Jvybs+3sIAus/pBQ+/3N6XEGEkTul2723mzg+sFAE
CdMiDIYSYHIiMjE9kucpkUszBIRmuv71+W3froHD5kv44APkxjIOHy0EU/xFb9hBKXc8VkaKG++4
WkAaRbWbIkiPmh5C3TLXusC+ecVIas/ngE/Zy6jYsOSnXuH59xcWQbj4p1clYVg4zbacvogJfdmn
KyImzaVYqS1zyLMTLHPSpHToUD9cTA+lfks5Ra7u/LPP7fTfgHhr7VUvvX21mDclowf51m6bUdZz
amR/1y0Ckq5vl30Vo53TxSleUnBdEDE3wAaG0O8UyQFTVMEe5RfcTGRfAbgcP0jMNqdDZpm2SHaD
zHpXiaf9IRMpfJy43E+hzlxvqIp0yhPwFu7Wn93ClgjbDHaGKpPjuVDKTsNFvIeXqdgFfCB+16kn
D8xQwoWmXXE8U6/U4IY9zRY/VWT07EgBVQb+efhkPjvpo8GWeVG431FhLnB+/ZlcGjt+XXn9GRm4
5f0K359D3SiujiTjMKCuo29RBGIYVFi0sMDvHRsw4thjjGSgaR7pPIILcx28fRtgwSTUfHi/qXwA
0I5nx4HVMpLOxxzVy+DBK8W9lmM4j7Fk/l2PnUdkNgq7C4KMcVTRc3kPLq+L2zxs8F0fuEEHFh1P
P8fXoVtO/5f1Ve7yenMyt9hG8D2UYx1T5e5Edr4ofOARl22rVhEaOKQgJHvbKz6cRyHmNtNf/2Kp
yBJugMBIyxAO9DT+XG4/hPfCBK/YhWH7UFtSpT6YHKdCBfgQmD266k/Cht+anHJHwIf2VcaEEH8s
hyFxYHPgXd8NI3FrHfjW30W9Io5Vfd04zJoOK+6ZoFpYnhj8flop0rB83Q8YUuwIACgjZMk7DlYC
64kE3Q/v+TLBnkWG4exBeGtEZOK9LqpPWde+kCGIhfc1BzAMPIpYtBlCrY4Ft+mWe66rvUUlXw7O
uCsgku8zL0j+SljBT9AaJ6lluCAKfzezLHuR7zB+DN0PzCPa+wZdrXHHI07TVTUN2X+RyYoTbY/n
uebMgpSWkdvqUvA210SZaVUZxUTQQ3LUnS4rJRXlY3Lk+VZP+O5XTFlloEdYxY0MujDnGUPl9EuN
/onXtIFfYRUx0d5AnferATNl7zcENgtFjvczQBzYDW+OjAS8YV86VtsciELLhU+VaXgpTp2dJbl2
jUx8o/gHDmSVyaxAJB6rrn77Tj5gtMk5A05Y+SMBDtNs1e3qQwC/2Z2wMwxxKhbnATGVa1p+KTRX
SyQr5mSt65SXawYeeIPM6W/GCBT4q/dWQ6Wsak7qCeRXK+T/W+fWggaM6J/nUw5ZaYhcovXDc1wQ
I1ZCYixE87Wa1qZz30CjMVBtXIOvrE15YGJdUrsgHJBiYLZFMOXhAQbJvTbxhqwRa7TgbLryoDUg
9ealKj3hzwmjh5LVF3r7fCxdtbK+TaXKQeVTCeLt0qHpXKKXlBBmkLMSmCs+UlpZcnmyxm5gK7UW
3jT4gJTXbwBMKowwWfYiWyOpWyqYn114HjFMssmNns5vDrGeaNP4N+PMenUlKRzR4oINWEq4B0iE
8XxT0SpGca2yAuH3HliSGRx1uCWRet1A0Yc3vEM9aytLa9mkadJueGHf7HUtyZHlctOrIYlBsoXd
sC4ym4mlg2PKDVosloJ6fU1A9KgFKw3p2f19f7/YcGsl9ge2ZbBZaL+rWKXNEIThrOX/pq2uO5jC
2PAGqvEKlyNbPEAYyh0V8ewvdVGPzcRrKQyBLGuWuZMfeYYkz+uVPqglSGYG3mPJwuUwOTAVciGK
mDf03nfR1v9OuYdnphgL/Uaq21875soclXxDt/6naT4xHJFjESjoUSnNqSQ5WVi3p4j7Ox1BuTKn
m2LUCKF4ksOmJcTrVW+5w0L6mdb+Aqb2UwJwtzdE0KQTHtK8R8gUN2gVVUEnXcgKwmlvNM0ccW/c
IYTFsWD4Sdg1rkz6yTgi+xNowcfEJbghVUxHUE1hSstOF7F6P5TqW35BOIeuADW7PzBlE2SHNUai
nhzolNCxpm/356uhtwivuPM6BWM7kV4EKY+rO57u292iPD3rw268n1We989sK9QoqNNdBep+3oNF
yaioPH+tC0JKj42LhegPpl0GSTewErmzbBrAEpxD0cOWK/Pu2nI498eBK9taO+DRarejDOKuJyhQ
+9reBXQhIgK39hs0vgEQYbcWOGnDwNNASvxE8u/aw5HfSsFnX41VElayhADx7G+9TCVfPyFnIOBA
N/GWRE9TVOmiPY87pa4WqOkV5WeXKV6wQqj7tXX0rA7M8QPstXLm1M2LZTAVo2o4LgzhNh1rbOpM
tAke59D/EHfuLrgR3jFavy55MXdflNxurPIPBGOxANPBROcQr4wV5/m7yUUf3xz5dSb8h79REYZK
PtmyqtPZxkgnjJU0R1hAU+CKOxvOjiJm9iNqKhFRt8gopNuzE8fXIrXxDJRn7WoN2rqD3afDtbik
lGZPpxq/e3S9/Z+IaAeFU1cevJz8zF96EunT7h0rPmKycWmjufhkP+2RvWGDX8WZe/rEy0Ts+ceW
atha9SZ2o/X1GfL4NrnS5Rq6jSF80TYfhvVlM0mjG84EVDFIzkNmtgTClPLyhmxf6KknSBL/60pp
XH4zcew8ZfF1euVfeeIf1Q4zIz8X7jIOGgHcEu847cJGC+2ttnfuuuuH5pFjPBu68TDwpaUcRn+v
d3jlmM8w15+LnjDYNObbeSSJTNEsc03rtY07zCCKR4NQ1RUClsa3DRugy1/x0pljRDljs6HaZzrS
kmJlyJFwVWlErpa27fr8FnTB4lLxtsQ2bIyETsW/IzjDB0crlwKMk0Ywr8sIV45kpGIP7mnra4U8
64NvdYTvNG0NecHMcVwsRi3I75SGizk6UJpVbRX5q+4E6Ko2dlf64mM8hgCSHxQXxrjT4qZ7DDvX
DqbWl/hXTOKVv2WslBZI+lXjsypiFifpNRKSMoM+AKsh0ryN+NtmLmKp11tzFkaGYxceMoiQL2wF
gcVizwG73XQCBh6tvEOnZXw9+vJ3t3T5gt8KS84O2EWxGXwMGl0YVtsQ7nUR+6TBjFqUpVp3c9po
1YAyZS0FhBkPb/CFRwzjof73GM4/rKOJ8BtkxKSaKK42guiVMb0UKtlg0gv9Hi6ZiHnA2XvUudzP
hgGxz7ntvJkVc/dvuM9zKccLZWVbZBHqsrwqnWCE1/1wVoFTuym0K4qKd7eD9YQBdTLXc0f+nImN
nRdDlieBz1tOvnbeWg7U7sNyAB7zhir/3D+UO6Ki3Or2iF9ejSXeyffiCwIu3d1DZ5UGzz5OPc6U
1CEYSC6mg5htP+QpWQ8OiCZqZRaEbRO1rFnf2GDfTqhOOUfxSC5qNX14E6rKl8sBHN93QIB5f9/L
oSUKqWB9t3gKmO2hniU7XBGEaMRTdEA/pBV/EhHioUyi6kNxlcuq7voPKvsF0gmjgre0eb+tOHc6
Qv8W4gC6KZ7AWS9L2FXK61ULxH68/jKCrEW/vu7kmQIZX88lUZeUtQcY0aHmPkzGQwwSfkNEyZDo
8S5l1QbEkt3xyeXg4Alb50PB7xnqkF8HOB2xnAG+ng27GYWTV8jOUxqUsD4QuJKur7RBKhbutaj2
f1cOuycDOTkBramL3GNrSKWPLUO5VgX4mUiALaKVZBV4M2TlRkm7mReuBcXO8+v545Y0SvseYqcB
fbTmK8Tneq9eob7tQ85lPUjedGXfWVjmUMVdS0hVBZOTdEVQ+WZQ9RbKl+4uSYIWLW0+f+qKxuRd
QonQXNqsw9CDYIdAUEcpkMjnphe6ZJ58XfBuPGa08qjPX/DmDrWho0s5gL+/pMzu6kjmGH/8tWAI
VLsDEyEg1fnq8jT2pBVDuUILGyWaTu9mYqHNGzXzgNM1Di2yOWOl+ADwIV/Ubbq0mSA5K5SdWsBa
ONDDNUiluDbnnzc/+wUeNKR3Ykn/pz3C4Y80FHvr+oQbrAZJ86hHrGPBK9XmjP6frJjJ4EdjOjwF
tXO01GKxSp4rqfQRbBlGShfrWntwnCzG6YKdmLJi6KNMP0DbKfQEtmruH0q9vA6bF9bdTiLzojBR
WiD+R7FcufR4cxDm/WD3R7Ev0eZYG/jd1FtR+EiDn3bjFDr5Ejam9EUMs7kDd+vnma7KpD+8cz54
h2p/EcLNmmQuPHvOTKyzH94ZVWxR2HLyjiY6uA6FMd5ZrD0sJGdlrGoWzFlST9UOOAF5cftCMPzz
L4rBgo+mEkmi7eW6iNG4iAFb1853ktgdnk/erZ2f0FVP0qkMbf1SqgD9R6UYc7CAMVKuHbB7LoUv
sCb7TxLJTsm4/JVNdv5TvcFOEYs73wYscbimyYkI3H0VjvBripxPbrLqFtW7+ifEtRvYXvVp4as0
v4tGcpD+Bs/edrZ923/LMfyuw2FsIHXZJR/ipsuEk5ghVZgK4VJf9bMkVfGRGcfAg0OfuQRe8vE4
sKn5rxmglTiv0udySxcW+1hy+7I1EiRPARVK7RkT4dqgxazXabzvq4ppyOMx5Lm+niguSaGX4eap
XW5LAfjumZN6DTYpnRAwnefHvgz1elUKSirdYCbv0ZHp6H0azFodKJLWKKobf/NGKE8gIgVJCxDM
pzsKqiZp131BCOZsU+WaUrQbZZ4fC8CNmEs2rbwUFxob54Ya28Rn2RIFoJGL+4AeU7v+OtZnZ/yv
otWhRZq6wQjSFiQrIs8HA76A3i7AdY1i/5jojdtj0/Ote3/Ri/5Ie7hPLzUQpAOujzq6XuvYeyYJ
5m+LXELuje7ZdobcL7d/bMXfY2JP9IUUqMk2m78rt9gatvbxyLQ9AWkC+rGdmEsJifEI7OC3Fd2k
fPwsekytzjC/YwAy/NJEZT5MxcgrUByeuxdcXdebzMsqzS90G7Oa0pOFFpYiwvzgLMVgiS8GLUDS
7qXkgXV+2aF6gwsQ8H4pAjdakKBIk80gfU5UYJk9p0VyH9AC4HGzroz4/OXni0Nj9uYs89KsyVeF
gQ+rjEsAuERdT7t4d5BWb8Rpb86iDehejO8YukH1P6DqOPFAPowEWck6vJVp1FzMKhwELKByT8St
Z8X9tVOwge+CLfIM3g7w4I+9gTxz9n+54sNoPLxcJu4WRWzzQCLf2B/lOk0+tLObPB8caGwWbpLs
G3LtE8ocy83ttr2WA+1jKac0Z67yrucVFRGgwO7ANyQXeelxLH18HIjrVQdyIFRZJ9yDkKKLZcgW
dTzzXUzfoJXNgfwDUPgcq9NNMpGMJsRlZyrgXZckFPFFzrgIJ8bzwWNPvG7ih6e7sWspTFcJsokE
LrrpAX6aduNZlJKQrchgM/GPTU1BYO+ghz//ySwKwEHkRRpr8v8ViJY/g28JCB4rZhBng3WG30NE
P5RkeQcGjEjeToptcJE8FLTWOF0CtCKMUhEysiM1DJ5ppI8wi910kGN4j9vzgQ1iQinZFRF+7+iX
0GPuo5B9F7STXjiQOSycCWjE15PoG6QmILPQlJQfj4yP2NHxbCnFSfQqJY89zNwf3NgEC3KUjuda
95VU9UnJ8bL0fA+c2fyfD/L0T7FUJyeAEF4WneFthyZVZC9vrQ8bcEHqyQ3EwBNC51nfZpn9GrpT
nAiBrg6OMi56Nw/QZMHgwGT1Nd2wJnklCvcMhRcj48LPIhj+pAu+xzTwM8x2QaHmT6cYwM+8Y2+y
I7u6CgpXt8FSkhf6y7BAd8/GZVJstHWuV6C0OaAGehLXJ5Qo1vf4kV7LhE+/Q3Y/5bOMXlolQ2Bh
I1OIGgejJCKiyj3lqxDih5LcfqJDIQ742R4/kJRx3+iAFo1vi9EWBZ+GoIVvkYzMg8nJj2guDTa7
+Cabzer8AMojxjoQgrD8W4O1IIbG3umNDnGf5Sh6yFySsesIFFRudgq8ZW68gjuQ71Vb4l4YKG9s
+vTy8bXcYTiThSbOdzlx/u9iIrL+6xXWcSxoa5Zcxuq0E8UTaI2k6XV5FpePL6P+92vFtK43xQ4S
0YRudrEmQbBxM5cXp8zp4rOTG9WI0mhmpTj91sYDfWB3VskJZWUfOBFFFEjuKm50pGiLIw/D9HCp
6y1apOl/nBGfgeEv4JQgm9w+VgaH2j8YVaJIosGqPqg/xQa9eNkDu4B+bH0TyhhSjc8Ax4qClafK
S9jqmXSfUgPl8aAb/0Yu66LgVmCyIHe821sLdo4QMEu6eZTgwbD4EK6Fyf8ksVukygfLm34OTqDd
Mmhzesf/MyVeDXFpyAwEHix0pelNwlpVjUy6N1IbNWzTvDBwzKs0eCC1UqcjwkxH2ZNmJJGJurmm
rg/AUeOgpE3CeTGcXigADW1gT+PTPx+NXon7kmtbRgOxtRr0Y7PiTlhrEJPtZseaMv7cj5jkwVg2
Xw7vKqnPjbFs+rFjwnJ1wT7vxu6FPJ7o4fk7t4wIQSRHc9GO8TGYiWAD1IXBkTy4aAzT7A1WLMxO
x6YIKPNK0mswNHaoTD3I/tbleeux1OvXZWqhxpKnHGPBX/gijRQArc2nMWiWH684sBznNWyyJHVO
wveyPKBh7iojt2hXz4nA+Y/gqk19qJsuRBClZCIxpGkhJNXmVXJQuyXysJDT2x/bRh1+xe0Em/m1
CW/t+OfKEwLWLUVsI3wFc1occmfyB+GEnGW/iehuCz5oLKY2SUJKFD0BPrx6p1imJQRpSdDEQXp1
QjRoze/S3b0J/3LG1HtRPfRor3B+mVQwH4Z8TEERSUGJbyFc92OTfnOJ6no2K6Cwpc5kOeAL6u6a
UXpb3jrEwarQuqjP01+7uGPFBEwixPAXbBUCQ4znuaclfeReSqH71aT34zJ/rX1lXznS38/FG/25
rWZACEVg0u2GcOQr/HDhJd0xQEeEqaw3X7KwCAzKMRxIegbXv8v+BRkQk83PaWyQIXVnezf2ij78
mtOBqOjA7FYX9zILsk38TXAG4Qwuj9thSRFdgJut+sKAXwx5JIi8qrFpAxEEbONTghkks5+C2QSl
P/VHHwHRv0/sRlz+5Vvtwb460tfhM+a/QFGq+f2rT8eS0kW1beQzU8k8fwQ2WQcpNV6m1i7VCfSq
BxKi8R8/IefQHEFa2xLwQqX9L36KKIcZU+/TiWlhZYVdtY7V64yWYzJftCL6E8bTRU8DtAbk4yHn
KpZ7ilZw3/7/X5es30AQmqDA3For0asM2nJKtu6p+r4l1SRFn1TK+VVPYkZ80gfAjh+pDpGFXrVl
Hlvh6WbTR1UPsj6IAUOlPcp4KMv0kKSPZKhydjgDV33XOIm7b8ibNc5BII1qbCKw08YEfQktokpO
8jXRNJSe0u/0xrniKHnaQG1AIydlaUbPN+X/6Ze+DHdeV2M7+8nomrazlu8Uv9/8wBW3EadHN/PO
TrPMRbZiMN+kb9rUimreX8NHHWBu5wCiHFK03xQNuwQOibDN2eZBwwmYhRavTHj09wDN/qVQH0GE
At54mRoHOtbwiRcvHWo08oilCFqx7TNPTOi/hv20J0a7qqNY9iqKMiyUSDvG6YQdTC/1PfRlSfqH
MxOVMJkw7ieZSHbPVgjq81F7yIlfuBUGUCDxHFAXNfq9Za3S1ekEuFagDShwPWu9cD84J5/afST7
hrxA8yScYckiF0IlChW//3oM9FesLSswkGjdQwtQB5hAdEcNOjDKHsU1XF3S2PUFx4Xf9pULpdET
WzHN+cELZm7+3DuBirfwfIE6LKIUBghP35LYSooLbXoocnTtJOLlKeZMuEODL2qN9jC+ZfCJ3uAA
+yBZZawkcfKCgi4o4puyy7GLatJBOY96AtV1n091x+xr+TZ29Y2EHeLC+h3BdMnig8iQkoldtqO+
Sg84y6G/lZJC1TjJ19OpiWsRWZ78tRaigQZEqJBjEEe+p/8Zoscq0ddSyvbSG4C7R35dW5whl1sS
z2kfizeDrBO1f+nBIwMizYgwKC5SiJ6FV5zd3I2jJjAxoskIjhlXWP0xOG6+DrXSi1zFy2WS/w+O
cRzsc408AM4BKTqJt3LCdPuqaUL/m/tXIjtzlJkoslUEg4idq+acf5DzuCvXTVYOFcO3l+ENbK3A
Bz1XQaecpMYHUD3U1BncOOWB2ElSkSODY+JA258fwOg6ob5WNHEwuGPyH56amluogramXuGqTbtm
/e5KP8Dyko9JyF/3M4T/zl+cWSm3asA1bxgswKOU1SdaBLtlpg9ydhABpu4L4jxv5Z1bd+PwjZmz
51tIYA+yHr9ny8hII1P+rCOguKTVOEQEIsDbthm2Kn1k0+G4TBStCWdoktUJMqRD5D8dz6Val3xC
iIPhEz1YPyRKMUMUl59jS7YkrRrEvGS2/+5SBRKe253BUVExrxpP62GE5mWs/2WGjaZihu9WPoFG
XOY77Aip8Ggw+J1KiN7YbTNms4tjtVTjbnOO9TGJj6GcvhlXN9zL3NJPaV/r08H9uwdW8brxAqzM
kga7VhdrE+Wo3DuSzn7I5AMgpWtOiRGSFhFWazMPh6ONpsaVXKTXi1Mp1CCIdxvmSR7fLsb1sOSU
iw/P01G6pWvnnUcFR6J4W7lp1c9yys5MrNowH9GP9zSrx+InnvNd8aJKqQ6unrkg1OWf4ybbTT98
Qi0zC79THgCrzU3P90swAo2s5G7SOhNheoi6psPtK6HlEJU2qVCo1g9/xo6H5Qf02757BHdZi0Ab
SOpAzto/I/izC7TJEnEGy7dNfjs7PdnWNMXbTqGUxTFwOnMsjKyQf/BGE0xIefxcREZg57HTtCc3
KvQqdrVo6zaGPVduL8k3mJB2pqRn5R3hcPJi4IcKYUWC6yO9ZFH8MxRNa0BLSy9+6PiV7jmjFRvR
HsFjr2Q5s6unUSKvyVtvnr+baINkUUdOnuzTqQ9v+gBnthCIxVY+VMpZRhnCniPTrDEXjSi0ERz/
Ot4Tk0WH+t4tJ2pIVmxHdlCBfuOdmT0Jy/BxJj+swXq11GMJGbfwtXSRvAYExB88ZGANsHasJz1H
lAii0p50sG8dI6TCSh8RTbxZK8Dv8zHa0mBPMDSPLDdB/5htFsxedhMsZAaCdOLdBEwp/j5BKetw
UTBfIqDHVhnqnKY3XANkjVKAhJt1Jlt/0iJ4fHcUB8+b6M+cufpe9McHBsfQmWiMIu5+Moz96MoA
IfkqyPppIpdxa1HKX4ZMxBj/XGqMYOKFJRuWptKTOhRRD+Qzw+sg/kyLvCYvC/AGVh5lzb6nE9ov
YHOvIR5ZDLW97K6HO1O7lO9BRo8nETTxuzK7yH81X+7dfyML+73ZvtAM9p8dUhRrW8ErR1FBiPF5
PNT9tRdMUQuwvK1wVgjOXkp7dddWi8IcAQYlca5B5iPeSTwBaEs0LlXCRdBxM9724KXbAcZ4Q8AZ
xxsDPD8El8QtPbE4SkeaJV+K0xuR3k8xI7TodTD4W3KNcOtWbPq7DXoxFuaZlDUDId0iTTxglFPB
d117mauDv3vmgoP3LsnxBCdmIw1OId40P4gBiOpRSjBy8Rb2lMIV1KIAup1gz/5rAiY2tLfhrL0d
GZfP+QOJNuB42G4LLiFRhjvDfJE/X5YQFLRrcFpGSoUcFgQZgF1iv6NRR6XzCJCbE9j5GSyvavA4
fngRaiZiJLnk6nBvXLctXrPxLsw4LNYL8TDD5AoUOaAmAnjjjgr7C8cIGyHnLn2Nw9hDXR0al26m
HDJxrcixprcWuqqBgFgf/qUzoiGVeC0+TmjCGWys/+ohfm28G4B9CeQ+A6fXy0iowpYi/LVVZ20c
jBKC4CQowl2OBcSSJUM9MK5HgX8v5PUJIUimRyzwgXsqjBcLKb8Od6RLtC16V72iter1D9VxE9uX
JoJEzvVmI8Mh3JOeoHC6dq9VE/IhOGdRJvDauWII6JQjw/FW3sNMFWWS3JmzLZ6gzQP/2WT4rjc5
obXmUzBhk1QZnmtxjVgglGpW3vP/EY6E3MhmvJ6i23GE59tfb3iaEOOvnP0F33jkUZMrMnnSVsbb
wHNLDYwzWNqcbIaSIdq0Mukx+farVX+6qp2cLmXBq3sKouj6aybxaWEex2M/8keNk+awRyAO3W/v
qJ/x/quWxEaeGoyN2Wjt7qSeieRV2M9cF7KdT72mMG2vNK4jImr0qC13P92OE5XvQctbhcOxeUe9
DMoJoRY+0Zq+YiA+31Xs9vEMVAYcA4TNaiWYzxR5qRpTKrx22lxU/ABFz5YAz7DezQEGewu+oA8g
eInQolVmM+mMCxHxQTOeHpXk0V4OMggBolOe6bUbxIhcnpYarjOCrh697zigzbcT+hBIh18W+hYn
uoT56GIOoXveHCvB3tc2ZMG54oFoBwOfsEBBkasRxhhTEPoeeaqwjTUeykOCLIn0cLSj7UgqdK5u
HOPIJ5jhG6fs+i6ygRaBej8UVqeZWy984Wd4ZEMgKdtxG9sVDXB2e98+51R4BpmbPofyjMU16fUm
4Z7ToGW8E/6OP1PyE2FBUXTuUlvixrJgKAjIVOS6ckQsLd8xLnfyS4fNvX72OKWWkLIPEKEOKxnW
rZJTY4bNq/2lxXVDwVJfgmODAn2cTKndlixB6sBMIhu9nj5N1LkRr0C6MvFKyzGEhv2dqvG6h6Gx
ArCnrKI1pdqZWjFn3gUwhNmRganPhYfX3Z5AhS/VOvrDBAknZfzDTS7XLPAjQOmixa3A6FbT2oTM
V6motA4OTvx9Jgja6vOqidt+cPLohu/0+4cLBgMO/f8hbFyCibcllFgmziwco7Y2gPl7j9teB01W
5nTbOUTGs4VpbpjCCruH+/oUV7M9xAv/lf9JJVjN7l+aOtLWn6+3cTMEDunUZ/bc37fMZG3TMEx9
4q4r68OK1vQUx2wO0HDMouvlu1pj7+Di6ZCL5/VmZO2ROhcG15wbyP0VmlPqoWoUaxGicn004CCN
VYtuleWBBaWxL3kIEF5QG9DytU02WwzhBq2yRfnDSB9pdFOINSq/r/n830ExLN0L1uuJcmdCIian
t/kt/e0DRcRpRk3h5+od1AVltmaU4emy3rA5PA9ova9LlUvI7Fz8uT+jTbys6byX0xa+OwGgcuYz
VzL+L5pmQgv3Saz/MmJqCAJK0rl/4kAp4GSz5Z1u4lPaLQuEmOiS+oGTSL/sR7ayqpQ6gOO+EyNb
t180jE9M6se9nKjg2rLucavZuEDmJGrzGGmv9JRNez9Y4lHWTPma1PgrnVrvJ5iAcy68kPlWOSCD
iEzyjaVbgEnhUNqVeFcpxisrqgo4EF7sNNEa5bIog/dw6gbfMWVP28O/CJYDFq6f3FzQ6c4ZQvMG
o2DE+ld+Ubu331D2UUk9BdX6MNu9yF0EGisjw2mMrvBp0PgiO0rQqyM08ie6gzooyffPJocYVPYh
IPEChMkf4ptBUV22suifF4kleRKjwSEviOK9U8ywGoXi/OEUOhWNxV8aPRcFXmWX7SX+1EItrHb+
9H2lJ8Qq5g/W4ZmdJ8lHzXjk9bASUaDs9L9ac3CV4CqEqpEm+TdxlrOl0PJQLPkLdboq3pb+dqUn
htJTfiKbyNDdSS/5KS1mlyW5pWszQVHun4e54Z6X0mfD5U7UsymrtGPupzT1o4sTqmy3F43azLyV
qYVNQ6m0oK+7RzdTebdkme+BOXO11xFQ16nDi1R+rZ9oeprYSyxZ4co5aiorBZ//T4+CUwXVhL4S
I2l2KncDROH/OxHILt5hqE98fKSnDr5y5BgWP72S8NaY58MatPTYd6ryRnakqf6m+jgMhR0cqddZ
QgBW164ceG17Yh6lOldNq2hx9IlQ69HSRw8aitPfcN9qD/TxzNXmHnAb1gnAyMRxlNm4BPFkQyME
zYhweclEeP+R2jyKRKpdk763QbTcuEF1S/AXz0tKwYclKB1N6/MciqOlziYhDY5aKYYLB1gueEVw
OFK2WOclicozTAX5pz6wGTVilenvKyL0OnaaGXj0Fg8qKsBEKusyga5f5n16n5oYqey4jZ4FJXaS
e+1/I7zUFsYMxy//3WO9o7GF4ZxmRatxGRWzllbUjNlWMI3LJGdm2DEIih1xHORx4S9pZAgnuoXB
+smlYhRERHqbqy7fsy+CQMzk0Vco2A923J2F1jI9V+qrl86IDs6Yn9vWgyNoBBKbY7ocKFLJiora
ZCCg75LNj/Djo4QJfxUn9B5Kfn4mOtVS6HwO4FeNKHcCdcNBjBmI6aUSmsGl1LbhHIRteo8Z/lH/
jbyIxlWztNqNWt8rp4dIHgq/CMOcB6096+klpYr1SLY+kmJrfhhvVFlZpi/lJG5QkRt2zE4wUdNQ
cJhA2IJKqDh7mSuaEmWS+OVp3GDARBvhhN02o46oWWzY9dwr/WxwKy+1zJnmiLtJ9iFwRKLhzuYZ
z3lnCDAhj061hi1PkbYJexm2ohJ4mar4sPKeK7V+D+ndtM2bs7qkdUL+klE0qaCRN+gHAgwGjS+c
sE5w+GPceY8FeuVRsr+ZSkVr5Crqnluf/UdiulceAdWnehGIRNXOQKZgUwqE+K1mmzxQZcPuNXAC
vrrZWCuVvj+/KYlOiiuJZTgcIFhhEEl1jjy2Q2J7DFHvjNZ1Cf2ntP3TuCLtX1Q8gS+OfanKwpkx
ALFnmHqoO0GV9MNHbZW1cd63HWixJvCjEtSm4FI4skvGhG5yTzt2CjMJsH78GJDf0lX5vSAstxih
HFrPbC10gHV1nI2zCNde5m9JCxcZAwz3fASgoF3cM8aZU3ePZMPJM4JcRjjUf3i3ysIv/9pW31eQ
yA91dNpyqxxCs+k7ws/FnMakKCMPBijLv6YU8X5ET89rRdrBInussGDUTgq0Fx5Uadvr7uJWPeWk
J97hpFZaZidyPI/obFsTMnF8F57Dduj3ntanUkDr7RZ8HXxze+5Un1itpsSDgm2DLexqfqIecc7p
G/D6QmLjzYJeLV+Cg8NviQoWOVdJ05k4Dq+0Z89o35z8+wisgh+gxe/PfULzT7fLls2p1Hd10RYG
Qot3VMxLdluh28NQQ/PEo9Zuzn9BBUWNlo7L11JXadsbUlkQGKYk9+3Cr9gEFwJZnBJnF0AMxars
BGHuTcVPclIht32iHhVRHDA4DoUxQixvdIqhrIymhOWkkg/v/UzH28motzKtt2WBqSPzlxgxW19I
QozFVuLB6NoflaHaYoa00/bYrgWwUX+YL3Fv6ljRrtX4HzoaYYzGWiCQZD8HwY6fZweN5x2i1nQz
wIovJC857a3ZyfVAgGcXxX9TRkk0ekrrEM4fUr5Z7P2Vp22pUaGbnslWjDB3M3DHMJpKS3jBjFVW
7I7kHJ2Ys665ROk0bUH440XUYmlofhQaHY2vT7CNoSkrjQRdj/R45oS2OjbtCZwIUG4RWJoPRJ2A
awSqolN0bk7vIUIgcXmsLUAqjwZxB4xfrDoSQQEE+ZoiUzkwapJxkZqsapt2rsLIqb/QYySar8a6
sJUnMAT83j8F3QJ9Ni7tzxedcHFSqSms1qufkTfK7iHLPnKjFS1po7DPmrzbsaD2Wr4gvYBHJh22
SIDqVIA7REflsjlcuY0oZWnu0IJK9ogEP8FkcC1zs9k/i59uhLC0mFq/VPwOO0UlTM6HxxcRvBpt
Y8am+7soTbbR84j3v2e/l1WQ+n48pWvYQTeK+qShTUBwcORSKCvVyRG6ZVYUVOVoxDpt8bpXZjhT
tRDXRZbV4jT8M41qW06creXjaI6lOaOEU62xyQkdqFvFiavt4r8CxCG3HqL3FXzBfDiXRYtBxFwP
jouMCKg49ClmzpYj6HF3sBBeVVxhOudPZGaGIRh0gstsKj1f9HBRaJz66CCfjoldiLERmjiNoKkS
tP0wuPCXj2wRxxjDwHhbBc8GV+G7ECVwuA/gWJubLuZdhMBaGw8uIjewIFJH7KS/JwKsazCUlzh0
vJMO9VkCb2tPR2t3pbh0HBQ/TEVW1FAA2rU5nyHK7Bok5raSMd9fk5Ja9Cn2Zg3qst+KB/frJrv/
F6ZolFgH2Euv6H3k4RWLtCHrTdEa9n4s9KoOd0dlubdlOFtXOnAA88hHQ/iSFctq0OzRa/UYYiYE
FSIBVJWU9pUZ/kc4EVE6OuWWVMP+kavCXicscyJp+fIVmdlfN2VXx9+Qi4ymerXpF503cFipqO1w
sRTZuWaCxGAu1t4U8lljqFSowYdQ6zgXL7dELIu3t93f+s+AgHb/NCDbo1qo98Kgob0+/I6dw1+d
hlNJFueMTaVqX9U5yg6vhQs41OW8WEyTJy8IsZgYaEDG0qmaReYjt8i/Mn1lsGjt89Ol3vrfP7uO
GettcHHwgwOm7AybeurvYixEUhe/0FcfsbGmruNcgXIqywxj5YoFnSgyD9BpwDKd3MjfNzmDmcL/
N2Dd0qmz+XUlpkkh4XlmeBDSN7xKbDdd23UMtSvOSR2vRwG2x5fy/1LfWB4pkmhN2vhoEC6h+2RE
bDPO1KMvOzKXmfrCC0ecivleXyZrc5IajL9HP/mWVBcnDEg8a2EWSMRYzu3m43OVlsPbpOWWFVJN
24Aw4qfK+xomVhjvcgKKIgdhoOI4wsX+lUhMc6Xr2WLSMD3YXsM6qT3ISOvzSwSaxMZ38POi0REH
vvwtSw6ngN9hLxzy4Iwk22Yn1EhlZmWzNm/bPkQqDYzPIONgDziXNuk9tg1MXXnezioFMmF2qzlH
gkb0wWwwgotMYOtKsUaR/q4gu/P2I6SCXUoKRYY5ilWY837o/+RgbDXAHpzMpKsghbKe/MG8bSq3
pYX+pj0noGbJpBeOgxwtbVNKJm1PRkjGN42cDBHUwhaVLYuw2yV46dUovhxeFsOpMApdoIPazulD
MTY2dZ4sxhN9TOlnZK5h6CHu0TNh9pqpXR6CcjZhOlmEIoAuNPr74c0w34egX+S3Gz6vF7cGQwnu
f2CiDy3alibA+h71SMu94GzasqqbH6iORBQRqKtkmXSm1AnCIg4s5WTDdvKYMVk5btLGo84Y9iK4
KTRYUMZ9ExJMFSJH54T+siW22NVPa6vZaqobVqP9AA9m+0SSw48TPNaST9yeFiC1zdtyABTpRxY9
hiFKSmVwePD2SMDRLY3k7Fd1FHtKv6mjSQUFK/P90MZIxDErFE68FEiExKqKGWIzD+Azoh18Obnt
hl3SglVjZhGiE6C7gwJ7sb4YvnPku3r+jeHc9ELJF6OuCNnLXaPFKcpKKmviryAkBGSSUYWVyuWk
92y052XJ/FiRD8wEOcPbS/uIOE8t21JTOn1dkOKx+/3heLZgItmhfNkE7hRudnOfDKAPyR9SOily
2asnZ4oPY3DkZ07m5DqLfgThVmNcGn+1Sp6fxc3Aes5DDZnynydACjiP/+ZU9zNiLZg69T0cb4yG
tDkvymkXFHKUU/u4FcKScUiThJmC2nj8wqePA+nfZUKFQx+3W0YWssHCec+Tu4k/+3dBoZazrNx9
gnVIgR4fkvIOwYhdbWUU0hpt78nHPWmtgCYQV3h1M9VFzYNdt6vzC/LrL0bQhnzu7hXb1oGk/cZL
sOkrsWu1w9P/88sN5mqfkk3RVU8t9of0+H39D56jm+JnFgNlqwJ3l6fRAQd4axEdQXrtwb8eth4g
M5AEMuQKZsbYuASiTUbVUA/Lm2TwzdrNEK1uT5yRGJbB/+dSIDwa5ty8c4EmTJFWXz2a/NCbi9JD
dShRt3mMAMZ96kjIWl2hfKLDt09NhRs8w46deVf6W5XtYBDoNPEZn0TA4Ohh1xT0QIp0lNJM6go6
3NacNXLmSRwjp7kt+9CGfICxsKXAi296WTt1oQGh1AMu+hxjYuF+xVHHtxpIqKUPlDeRnxW7Dea9
8C+7VjywsOsfv8+/AjrVo9tKhDXDXj8JLQDilGRDfiXThijFuGJp3SUjRK9ZtGPNpfHpSnrHNewC
K1mxjFJoxydStjdmr90n+MbzkLjJrhOlIj6+/h/j8zLTzUIhtz5rRyIELinZAheQyIqZQW8IXv5N
1zQHjf07HN8Q2jdzLhVbEIby1kN4cwun+4n7Ubx23kd3Yg9n7A8MRUTbfYOuqq5C8cSFq1MhZJ48
Lb1ZmMtMu68X0+yXzQxhU2eA1zHaRTT1Ok4Pua08N+7b0I6dzUjfHN3juOJ80iOb3rvqh72zJNUp
cfbODdMUngefWb/Ts7YMAqQA/ZasUqnVxOzJ8pfDq5xk1vZuAgSXQSyIFsGUBZUIFaNuxzQnNV1/
h9OEGf4rHdd2kIwhtreQ/YojlabdAMJW9v3Tw0wjgK2icthhpCMmVDmR4LGxk3xnHfqMaX07XKwl
s2dJW1tCbsPHMd/Vo5Braz5rZYpCY48t97vb4Je8kG1SW9gAr88wilTO9o0xbIdDzQVlSj+36rWS
UBqbC6lmH/ULKiBkfLxNuStZqBF5p17n/6Lbs0R0t3jHO1KjUauGruUjVt730Qbzbvy7wobKm72t
pVNYT3RkBHeSux1WOoaujMeQPAxiBmhoMP0xcAixCOPsvTK9czwd/Wi6izxQUEeigbZ0GLY2KENM
x1b0DBjncu9hxLPOeI1wukEEeb5CdHEqT9O+OIt4DyVkOzdHOjdQ1u9kkJaPhupyz15vXoveZMyD
RDNOKb4bs3+dWdiaNQmr9ZaUvbhx9VOjeoUHTSYOPGjY0VFOznm+jb3fgWe52m5GZ2+vlOJ6740E
U8P9cJsk+WVUnYixYOhRcyp8fIQf9zP782eah3gI/qrNjmFBZ08Pt5NZgMqDyPNO5HkFYoamgVPC
cGYHrsMn3tYtoa+i2y5EAGUv/V4iHqu+stDYv4f+DkiCDu+gwnnNB2LJHVA89Ce+G4fqnzZa5MVz
Igj2/fM6NSVTAwhJFwS2ySPj1TIJpvt278hxCvFjRlnf/2dbwk3dj+7rw75O/4KrT/p246IbgBBt
pV1eFowXzim5O/u43XD4SKrdk8wz9Qt6Kfwo9SkNGA9p+bSxyYcFGQpBl64yHgFmpaYyodb653FW
gQpMjBkOS336MXqtSZtOxcL1SAfUXe8iKlpfWjRG4q33izWbaoX/A5xoIXMps9bJy041zQpPkaQn
XReAuasF9TF+GAdxKa1XupMMs2/gPepMh1ZXW8Tfe95L/anIEKijXbau38hti7vMs0AfsdNJeQnM
J9PMyuaJgPKbJJTWO8bqKxDzwF/qZ5BsSLlviBOTUbszS6lBRz4XwKkVOcOFl3/X2vQeihcF1FGO
mAmA4MSMA9shtUtWLY91CxqCLDhuYOk2ysduhyUz+KGGMYYjJ9RZ0Yq9Zm2CCN9ePn6xdMs8b4Ka
9xHX/GQ1sK6jyFfxwP8T84f/R0dPKxyNW9WANyO0+3lbiwmd7oePfMc2VbNYgypIh7oKe98BHwGy
RunfQFajR9zJQbdRF2XP4cxl+ShyunZcwmxUoW5o7M/P83egTyZk3UzRdR01xWJt7YkCbErfhrxy
k7pj3Gi7usarnkuzg4gM/s5BOFD6Q0N23J2ocN7jl0fOdnSov/id2Lmtevx53TTGBDK8mx5Nfjal
G2no4bXdk2Nshfa5k3L1JnxBuYyZ9y/5Gc2rk0wnuBuupzo5dfmVIb2oVfMeWKwZn4OPoyEu1gEs
mVZCwCOwnML/mr/ZpVG6+gTiGOmnne/GSzCuesJVny1tNZinRBjYIlcdoqT3Kaf+NZCP95ld8Lof
IqrFXga/9lBsqdXcVTzgBzPxwHVhJfZHXy1RHwxgUYwErZXNJv/VWXohN/Z5BqXSqRHdzntBCipI
UuA5EVF1VUJ+V6xQOzoPaDjph98Udbunr4K5qdm4rV4afqOZ2IIWmjOEplaTcHFSIy30CHrxJ+y1
eWtliguzo6rnGJ0ac3EZgkOWHEZofxnbtpLMAGrk/vrebxiSdCXZ8xS05OCJ9UyUkDwBmMk8J4+i
EZQ23pvLBE6zLcu5/kkSiYfTQKK+hPZmLo89d555laRQHkxNIrBlb15Af2Y/TbrDRW7Z+JCbC4hu
7ryD5VWcESORN4eFdwXIlYPt2o5VAPjW8hq0QjjidCTMzkTDVe1XtzCWck/S/V42eyQ4I4PXViDv
jvg66m6Piwe2iI9VQJt/wHyFiLHUXiP7oGUm33RGrMdyhIPyfHEeOm9UN7md3EkWeLDQkIyOYsK4
W159bZ0xAOKmvYx0LLtcYzF/OsmOBv0NvQMCNx0Rih7TloHE8mmUSHrDpNXBHp/doN0u05udx6Un
g3F6fvr8Tk7XE2W2juitVU0X+rBWT0wmIZw28/LVg/XDagSS9iBjEvPoHmjS27UzV1m/DrdgnSVi
tgsR7UvQdbIA7oV5VBdBmYEUEhekYyHS8ABswtGcCxQY6CG523eOdXzU8ltyxNJKOsMXQ6wk1o4i
yAbeBRkHhHgz5OSLgkJHTT3ENot00V4mbvaBRak7m3D2zd26w0Z7lPDDsslCli3RocOL0XZ9lq5x
esySbAATS7qWHyBeT2+Wgma/uCNxLBty1eSIHp67EmZq/r3k988MHrxNLgJLB8G0NkyHRxGudAH0
DfXrdzm0j+2qss1utKEZjhFtti7IBeqFcAAI12Mtox2k9J7Ljqkc+K6t67cXCqct4gY8IAo6HvNf
dIWq8e8zXh67Yk/Li956m9ZLS2VIcCcVMZkuRpfQlIX331nU4S7ui9FNRXxt4fHbKPIHBFpn6w3L
W2zT2XwDA8rjF5AD27FVAyW70LO8JE06UgcxDuGkQ6RDBHJqHJAUseV/LfLcmXDuXsCDUTD/q35Z
cE/MSAMlMwtcAICDoSI6PTZFkGte7rocq7erDtZdiy6WIOx0F0llON6K0s5eFxuycW8DRbjqBC+A
/Np8afinPTWhhVgo2eoP73bRanMHzbtn+9wB11sd6rWXP+oCcUWG9S+aA7NEuGFoi/+G2Ayg//M9
RBmN1qm4i6XkLpRas/YAK8n/aBIop5yk3Naz8WBHpr318f9TJoJ3DshELZkMzsmAiXvzESXRpYYd
bJwCey7TqW4sVcFBg7TfnDeC0XjptLnTv8FMktykHgYjYlfw/s2kYwhLBqt1GfrSuBRRck2fBgCF
ugJLwqpNzHkXOMi+DtcjwT8tji2UCqFIh4XIBnetNGInJot6JUkwaSi1cgLtbLOgO31NB5Y9eJa3
tGH3UW0UGL25IM5+wb5GFmn0bK63xGidicT9RHiQUtHvsKg0u1XgORD+zp/sA8RAn1TuBasp0h0q
FTZFY41PgFxFs2lNAGh2YO3JDY0SCmQFzh5rv0sOAQMEuXkWuH9avPong0k5hlqtAVz7vhAsFC84
O71dg87g6eun6Hm9h2Di+ee7ga7RZ4bzWzjM8zrUiwoa7xTACPTI6LSymIalMkB0lPhgM9yl0Otd
A+qdv8bhoxb7AFcpniT+PfHS+yjWTmu1kITFDLd1r2PMDOaLjaKmaObWTrGxp1rIs6ryJG5AB8Lx
Cn0P0RrbFU9kXKGjPHTWS/jegdLJMGl4RsdaGJS+v9SKritEt6oxG9q7LNGQOEFPw3gX2Lg/0GcP
mern2aIAQmz6JF48vgen0tid0P/pJAyxgUXeIjWcMPNRpkqZDyEPpQ9SPSqcdLhnFXLxfY2cC9Qe
BB58VVucFostX9DxYpLPRVUfEHnqsxj/eS0TCsru2Nzv11IOioE6fE2l8IYnCSMyOdJNhlZWeMf1
i3Nc7wJNPtl1WaKQQnwjm0eiZCNE06UvRkdnoTGlt5oLA68yDCVG1bgq3aVxJOe/d6OLCC/ONXSJ
NndXkTwWI/7Ve+raOWTUzYsbfssoiv/1YWnRDJ4twWzzwtA2uIyf+fvLx2Ip3YMFT4QBAI7soP9o
gQzwjngAnVR8YEomFgX26MetP9YM7cmHHVJWuVj6sg/7izYNPmm0quOyNiye14Qm9fl7nxQVwoai
zqTXl9eUqQo2ZE1oa/N/wXPJw3Yj5xAerPFRY1wXXjzFV6w1Phz0Y0XL1of52gvABDv4ls8aBWfB
K8hb5Lm8ITJPISe3mjlfEVFtHL/VVSWceYfqzQUWkzV/laYo+0z5AomXojunT86y0QHuP2dRRZpQ
e0QB7PkT8dC6kT2uLS/tlVU0RnZn4sBDt1uWn1ctOXgmgUrHiOwngE+w8vRZBtSIIArn2HY7TEJq
Doia8pdrk4Sk5Ihmf6B3OeN/HaiDnM4ptTeu/BV8cEcqKwUtHD5STF0mHLgmpjEgjjh7BD5FKLGQ
uX7adfJ+7ZCr6cVOog2xtUU4CPz1odsmICveBJTzIsPBwKhymi3lDCJ1lOeB9pI782fYyzlYwSyT
hr30ltlTFgVNAAAzSbTUmkBvQlchpTfKwI7wfHF2FVWKyAJs1yrZFlhjYgSTU9W11IBsfB6QJjsZ
u5fuBGMClScKsRSAyC74HzdYPsUVSH3Vn4BCWVuq0XffuugqdM+QKk+WIBtrOxSNdYp1D1ZCZp0I
S7WRJwZVkYAvKd/6FkCYi6+0SSVwuEpS26hD5NaQkKE9A1F6upxa0SSTRiAy4QUSkpExtcXiE2tk
kJ16PrXmp29mIIf4Mjv3+onBp/wrmeDuOFQtw8zJRhyYdZQPB1t6SuhvvsRNiUcZ2VR7r9MiiKiu
TYsI9+j7Z0q5l0hNd+KyFIufBmnziM0oC6HQQ8aRJoHGzZ6T/NK6xXY8sVxRvmZVUKV6JK7Q0T58
ADWyH1g9RPDnvd6oAxurfUEE1HxLC6UoevbFIkDLDdricP1zWSHGP2YESZF1NLi04M1kax+5ofNL
9KJxxT7HcxbnIhS58y571sTRKdAlFZsLkvBRhO8XUzAhSZVhWOcYFsO77VDvfieHQZ5rRHDNZuXS
h2JPTIX7ibqoMATkmHjK2F7lwXQy1XI/GB0cayS/r6xQlcOsf1pLFaKzSIbqPL8KoWU7mqXfk1Vs
j/UQvGp3pEhEHpbv8Rcg0TEY9l3gViyGRRFFWZL4LJ7NiGGyhRNs4onx+84mgTywdADjQ225732q
TEv5RrsyH360sb9XdTgL9sPnnWlwVRlYSgFH4rblHlCQsAOSyI2LJD7v4XSaynOpJhg/dLfymug9
hvnF3NCvIxIdjAeN44dOHSMXWJRghpj7P/d6h/qv2FFU7AqcZqK0XBQ9PyqHipvXwUYgv6QR6NLk
WMdTHX7zDI1X6p6QpcP4mjozgVjtlrQZC1ZGM5gIRoaj+sB4RZ610OVeoPG+nHIutIljuvhmCHZN
y6seCYtA1KzZUdaa2hEQcB+5k4vV6tOFEmqLVsbsfaDtjmaQLG+JPE9N+KDFdyBS/6nCtu9J3Z9O
LT/RRYWLupdJyo4fAuizYGPePcdC+AyB4v8as58Lea+UYZ6lHa01QoFfAVB924wMFLUZvIegE3J7
JBHO1CeX42qljFl+feeFW+rVqV3loSFRAiYGzWCXoo93Dtf1HfLzXs6hOgPbpkx5zFH5h1JMKVn/
LCJfpEGHuJzd3e+vWX9qw0H8VfSEWGhr9zvDUHpXyQI3P3On+sAb2s23ciSBS2rrDGqyQzgf6u69
DUiDC2enO+K6JAgI8CxznbBJt4JJBT+p7W+7Aq+vA6BONt0YOyTskLxTH4cu/uafckvy0nPUQAns
EX3uJ0g2bUagpeeb5ZjAJ1pbG1hDP+JgDNaTYhvInBvgE9C08YWl6+TBVzNQHRP+GegspcWV8mBf
/yVd7BRk12hbLuzepbhbbd5p9sOutGsu9uVCgYRNYc0eFfVuA/NUyY6FiX5vlyshI3AQquoq1DR8
afgZV6NvYEvex2s91fIFSEJ73tBXbVP7YogYwOZOImkRwTLFvDcd64UNY05LPW3Av+l/Ztv2E/KP
T3/edsVv3dYAfD3SbdkUp4XrG6PTVgZm7/Ezgy6WXKp4SkXxEqT9wwtrzYiZAY37ptOhOwcg+2eC
Wq4a2repIelXFBX82Fl4LKzZ/uCn91eEagX1nGb/Dnn1Qo8qWdEdX4GS4iUyCTwbMBLQ2TxzDxUM
PPQsYN+SkmQDQsGBLY+XGBVSpirIye6ffDivAbVqqE7U2nrqrNKvDpcyzHdc8HI+FXdsiL0auESV
1oXJwHuiG2VUA00J8fcDw937qYh2Z+AlmrRe6gaq15G64dN9oQk86s+2VNyuUOJEBBkJx1BSGE4f
DNAgbkByUgGftYIKuX6gLtM8KF9j9o3JFb8np/P5U4uaiMKSq3FAsWp63DVN+YmNHXUoGku/2KBh
jpbpycxory3VEOqpkEA87eHftsxVmzQ5cxoOAYDKeXDYUUKHC/YkI8SoHW119yIA01ZL+qg0x3mX
qFaIVgYOsvQSwjmTuTS5M4AqBepojYIhVFS5KZk6KwdQdAk7ff1i1I7pxgRTHSNHID8OFEcgjJIn
xST843xecgkj2qa4dJnVEmqL0JAasltvMamNMZnLRWOyv1HGh/VzghKbgfn6xdBODwYxPhl8e4BS
+wJshgaoqCYNVQSB4tr00wjS3g/GzZVd98XEV9N2asnH3QOG3Uhp8cUVkTzZwKBzTjvpp4S+0K1x
NlS0IsKd/YnzJ+/YZ7uT+L/CP9M0/cfUizWva+wap2ya3ib7C7WiFwiWMnlIX4ly9Smeo45saeKA
PxL8dBovAFTbswVGdRaDyTuj9o7TQErBwFCbkaU0eo7o/12VSTHWj/5ptCyLlRXvgIDjRVLzLLMH
aG6OsaUGTQXvPGnxe9JHFgAg9S+3dX8UFrOVtOWOIUPQdJsU2RqZz+qw0bdx1Bkr3vN9oijudARl
1EWdUJSp9zmk7Ni119jG3Gv+1GXdka578KmZicyJj1oTrHk61IGjBlbwKuJZnQkSd6JR/WffRETy
Cku9JROW7ng6pCAMJzOTfviMHoqRZdUUv46mbP38BgBEjR2kpXk2RODTrldJpDMqbejHTVsnpYbu
tfzb3lfmGxg2/4R7Yek2vMQj4fcJrb+Af8p3rjXnXV6ebnWqql2UXmdQXYSlZi/4ehawDb9qoggn
YoGECCf9F0yPXPWAb7UFilums+5x20EhPh1m0GbUWu+TyCPPBQkK86gGtawrIQISih8NfZgkQnBL
HQd00GuMsq8QrvHOjxfbp0mHztm64JgQf6dzZXwtpagkVMsHD80h31qoqsNvcyKJa7AUJNCixaOm
/Hv2MlVqAusBgZTHvxfJUJkCUkaIXZAgwa/14GZZLaQmKZ4KIFeIKMWhyG/Z4f/iYTMKM3BT8Whr
qTaAwNcoyAdbE2vm36klDwPsac7ylIb00MUeo1X/LLFwrpZFb6L4cd9lTU3WNhzcrERBOPLo0gK+
0FRvHbc7F7wr4Dzdkytb5/N0Fi6Rq72mKVqjBs1JWm5SwAWxwYzgNMvvhQe12l/LWQdfxcl34J/u
yUfkfSJJ4hlwfe2ZrJdUfFcuN8gNhTUPlq8G/3iT0yudSUt+foytriGgFmar43/CLvVPbFCq9SGq
kxKK/FVUrh5dh1iOeMRffjIqZLilwn6fd7SzQeyNPIrjHOLjpwHHS9Q1McoJiYl05TWEnkVpYmI1
3LBGpkN0QlciGlxEzczolQtfBMmorF1ridKj7cu+JrAF8MpdHOAE7/e03R98H3odh5KK9FKOnQbb
PYKBuiR0W0cNyusY5Q/jrvL6LL10dTEgYiU51X0W1Ed2nD3PP7KkXy2RfaDEFgZpKLdNz+qym/KZ
VLZexixYByjX7B6VwFq4k+zVzeQlSdNXP+t5ccolo8pXEr04SDV1ZQ2MYeYffJM6GHNQvGDOKuDN
4WD4IzSlTnM1q7HpQ7FhBSX/rKas+THOXfaPYIRJfJlWqjEN1a6kjLMROT74FKW2DkbsKp1IYJew
jKWUi+cLPbejdmrepGGl0W67kT9lrHkA/FqqgyWJtigarLuwWya/Vsv7MAIf+TZBQbFeM1ba2PxY
z3QgQhNxvgkukOvFl7ehGfWPcLZw9w8DNp9Ee0pNc2vU5Qn23ZnnDJN1Nkk3IooXxvIF4lT8bhw8
9LYtJ6/a4rhTeqiaEwWJIlJvT92bBwEEdUdYaEOnbCXlfni7hcdQ6hqqpVcaJxATBVRh5mCSApSE
04z2mURHAfz1fAxzlFMyWH/twIxxbDcmG7zT1wj/Wj5w2F+FTgxXEDPn8KUyc5kXVDUPDBMdbrot
QOlmQr48/Mt3vV03/OphnaA6bPYPK2Bo+9BvToo0Em0F48UgqjjQUBv74Fm9JrmeZ5P30xH98qjI
gXwkJmSagwpArJptoMTp76bn6WuJLKb9HPef4q//A/dITW1YI3YtAFQM4uUox8PjY3sPyxkzrjKB
QIEOAmWBCbA6OsWjq6ioM1t5zfZxkb8JvHnfwrzZ6f6CwZoS/fap+Xv+6ek7tWpvr2sstQGOX/TU
WMEWRvZifOXdsEHN307fynosapvfedDBfRLz8ecFFaW37uCdbBJG96f0dqPjT/V5nHoPNx0BcVZ3
1RKCT2ZKomWAq01PTkrdq1pISB0RvcIIztG5s2W8P5jDNjqgNd+eEDo+iEJapPY+DkPjHsjLdNi+
nGeTcWF4BlPXhcqThsAer7C+uSgZ1Aqh53EeEHk7GDVYR3ho905inAEEyXUXmoCkb16cxnXgL3nh
eb7DTw6dVrtPTWJOhRBKyJrTyOxT4MPoLdFlP3qymVBOPm5IpoVXZcpep6SyE6ZpPH/frD+DQUsx
iTv97nLokGv9pw3RODwqKbQ3igkB1vyfZOiCvmAmqMiwZg3p5Gsz8u+oe+EfWgona4/1pngRO5Qr
Dn56V43V963rzYKVVxv2x9JhphwlXCzHnIuL44Tbtdj6MBIuresTDy0CEGZ/OxcxO3WDEtK9hiAH
Jc5CKdbeurRJ0+EVI/zSOXvN047xBN6s8NrfsyHB0moaKJ8tKqVekM9pe3uXcF0sKSy3ulGFM7+F
GyQTu0bdbPrEq3qA62JyHr37fbYvrMUMXF9kSjnMdBpFJTY/PoA7ALuHVeEs6DB7ruFLgMHBsfG0
cANl2799oC5ocGTzKwR61V/qaj2Drd3Tv/lmVW9ZwgN7nq1atPSkM4LI6oO8OSlJEHm80wHJjA/B
lCOl3kh0SA8WEhAvwcJZZvLOQvFn2sRviUYPjVvDeGdT0+CTd3oMRtbJ2JEQSOyNYkeKmzZgX7qp
EJyP2CUL6HS94BSyQDeZShkUjI8om84+Iunl2tvzg0IS1l6eLdFngTESBR4qvwc1NJ2Rv0cg+4AU
9a4cm5B9hvO79YjX38r5HBOmldi+1z0Ujld7UE+qOm+XUYPfHh40s31yjVgtwmlHG5NYYfpriv8J
jzi6LZnr4fNukL0IrGhu19UzQ3kGZCIkejDCiT/NpiCZkKy6/KvpiBJwXX4S/22AYN/GOlUkXSh3
gOjfWSUSAZft5FaD2tpdPaqvJf/JcwSnBvyG73OLcTTnjsVCHEyMNSbEXjAg3I8YlLaaBrnMH65q
V5hmTybiO090ULPjprZz5VgPYz2zMhsK7h9owpv0WaD2nfD7XwYOny/n/VWNj4gNohLKNHLhnkG3
5qGhGUyjZR+i2WwR0A+2MB7IbeOMVtcb5x4DZ1luz/u/9oIaKr1u/tLwc/G13v/EnkbAk0qHR7Ov
EKTQp5hDfGFiBJYkDF1Jn9Xv/0oXXf9qOkpo1+WR3wy98DuT17zD8I+Ark8o355KH2TTpxHSEz3S
x3gNPDyMXgCLRHAZQqRGYsNylLXdH0a7pHWgsAcAOQRggCIxum0RHlvrC3o1mRCyrqYXqHmldPv6
wrjEJItvezdHA5HdSdmsAixDegVMCLf9ervOgzbi3oRGUWMmfGTqIhwBAhj1mwMknId5IpgF1Dle
m7kMhYLUcKe2kcqB8nZPmRHdlHWhS5NmSnPKnGxHtwW90kY2Zi2tKzVFlMArmi3vrMyYFDk93V/I
nkN1FMrqbaurPS9ItcUfNDrgBtGUUKV95S0q6oXMzCsLjsPghRrJsFOo1GSv7SN5eIr2n7bzdYM5
OJQOYDqZQL+Av9gAyVHjpLzhiXV/rdF8Ccdi0VCCzt/C4ObYHoGLQKPREbUG5DFYxFOm4Deq9Z9H
bzWt9w/LoL8gmWDwpgNB6/Kfto9MiQWna4evOgxVaSpt4ZIykxe3JD0iO16Tcaj7NPguOfKeyr0E
wnRKefKoq89CAlSfOF0WihoZkLVEL2g7zxKDbfe+Bp+yg/2MK7rOyPOBUFCnIvpJ+YMVZa5o7voB
5ww9sU6Hhn9o+rWWChdP0AGy16Tr1k8XczaB4/oKNVSRs4HiRmRQ4x4RyNkRo+v9f5x1iyzRfQYI
Nr/c83+JY0fW0kFdRu6Y6U9fiiw7FAsCuOQl8tupnGbkOk5Aizh2uCrH2zK5dv27br24V7PxFGNn
jPxolQzG1s+1bvH5iZ+AXChyuynupCkvhyhPboSe1bOFf6F7HnWvLtSX4Hf240o6hRY3+AosoCfH
xzXEkzAyPjx8BqFL7NBqiabxPDP5uOky2XK/awv67v+69eXNwMOWS58HnsHYWTbGnqoTSrV3ZX5J
Nt9SSSKgawpWeiuGIwRBsmWf0t1LsoWw1m9OPpChww+d4sHiUjYN2wtM6ZyFmhT0GM7ZcoYsMoij
IgS+4XzgykhTB+Pel/eamlI0Ng1oiIVRTVoNo3dZ5+YXxLEB/YHxLLA0+FTln3UeGX6E9DGG1E3p
+8M8NCdZE9rUVXSQrt+gXvRmCY6Vm6uzz2WYOeeKMBht9CuCyNNQSv7KgvIS3rJA/mnFKR6aCf0F
P/+4yTG1P1GUzS3wsoemxQ144KkqkottNWZnhnXrrtOsiDp6xItbQZ08kRnyAjDmMdGQ/75GoL1X
FeHThCZsmCp0TrtkRi78Uf23xKm+EDfgrIkF82FSDj57YZM3rLfGYooiQlHMpegf0gfT7P5rlI2k
zB73U/OOf5yNJTjlbXy23GsI5RdJEcNsiiSArfOrePVViUR5f/XlDkXCVKRc61mwlQz3ue6dNy/w
9nWTQb2FYIaZ0UihYIre06KolYAMUBIqe0HClINqK1JdctB2gSDNPQsskUkevfuzDSSx/zJQbRBA
A+e0/AAubCuXgQfuCGDVAB6rpqIC34aLvplG28pAKTVE+EN79qGhNyf67NqjMuTJ8+SHKAPjqrG0
Nf5mQjaDfRjZtbNlNbUlcHnO/GoaQpMu73q/nUfHp6PN49OH1Lq80N6ZPEUjrdniWcnzKsRbilEz
G3kqM+ptWLO7XGld6+yEKiUeXvf9d8S6XOQpa7K3lgQFtiPtsNWXBHO6YVw99+U735nl0+yXe0rL
8faj8NhMvR4BrbTbsf9IOu79sWajp9hkAxlbWgQnOZjJXtDd76XKMsGG36RaKbCmDe1v52X9+WTO
12IR9FC3YdEKa/xWL9cmvV3P8kz6Hsb/MA4Mf+3CGvR4V7QUAKxiKXmNN+neUcYiI5iRLYSfFoD6
3u2vtXDwnqbHB8Hr/RqyxbPEQdvI8x9tf0t8pNt13/sAzIdnrd/LYg7M7fhzQL7w980b365tjGTv
mLfRcf0K17p7kZ02Mc6SB14Yw5m+HpefGFwQWu6ZxWWxF3M2dZYSNAvy937hqwLvGSJTv4v6GJCM
3Qr/1zpA1Vz4e7jQaKhpT9yW9HqUf72ivx5QQxdE2Q7ynjQ3/33fHTy9KAARXGmjhGK4LzdBMsAW
pEFFwEy8WYJr5LVYVYQONmNAaGsiKTEgrOQoy3m2L1/Nq0qZOofPgVWQycpyjmniq13WSNC5poeQ
KDSChykIHVNLAzFe3Mqgs5BiDEBH5lKJyc17A18Z4cX0VjwV2jd9RDucTzaXksZmOXSIXifk1/U0
vWZCehjgJQP9pVHKMDj9rQFH2UGpUOFVGLjgGSDPjSG4lTkw29F57CGnhRbAeRItudoU9ojM3jCf
mo2sqMTFsgYBCxJRQp7scBYSSGkF36mZ0EMoXBN8zEoHFmsGiNRG+EHzj0v3dZ0uIO+utHGAb3cM
DQYIk1Sf5BYpMDM7iWdrFSinP7wFQ31dzX8yinu+TfZ/ztTLSsfqgfakXTBWzCnZKS/0yoDpCD+7
KpN/AiwH22LlxR6HrJvmCLc5JzFeQv7Speqaq4U5+x713BHzCFmLOmv+BK/gySZeZK96M39pPtS9
FhkyeJN57EwkGcPwUXLQwoiNq1CHImD626wDHLUGGbLCFGEUkcLMu5dVGyMSMgSKa7fTCF6qtK6g
jKl43g9G9ZVCz74Swh0YAF6SUWJr+KCgi8YrycZmFHsEAg5KHAYTDpUSE3kHZtAbB4FFM+u58jr1
GkXE74F3NzwOBg1x35Uis2GQmcEnxxHsrUw8Q/xtfvPTli5BwZQpOmREe3u6zbsMr0dUCnnELrGg
APLKVWXdGwurEd8emliWhfshXhgP/O1APNH4pQbSMTSCjo1Ch5FEOoETFLqJGWyY25rJ2TvGLBp2
G9lrquiRKIa2Los6f3emxwwKtoI9d01KOCvvsvuhFJweOWiCbFYR6Nts3tiq5JBehJHy6yi2ZCUz
JPHm2GcoMEbjGfnGLwuccZ8kQCAz/jgmIFXaRoFC8TGSB1BD3TMr0Bep3vIO+XI7DGEbh1WO72q2
J4qmfC3/fj1I2KFmSyNLTapybSycqsvzR3r8r9SFtPFGCEFcW5xz4DgdTuJo6dDFRouIZlM0IPeo
vXxgS6F78BLKsDeC/blzqsFNUPn7pfKlPLwiaEED0EXq4Y/fZZposJjVvn3vy7YcHjJt7pWFJPnr
PmjO4UXCEBHmn09HxoEcHtUmKEboy9iM4JJfdzPt1/ScsB09M+IYgioHqS41Q25MYZVI3BEFKzrn
8I8O9UustIcR+l+Gvm/jRUcuJE/+xZY/jVHEkEo8YmoQIh7M2y7f9WvjBq86rK6/uMJ/2svHO4fy
SBXuSLj9JnCysU23Zq+7lGxBf63EU0f/mvioxKFJhnWiV0XoVpGb0V8S4XQZEIYtS6kb50BLDECa
Ty/rwNjvR2IAarOQRFVOW6Por1KL3FrLqnnDryDU4SQIGqDzJucGBGJMCbxD6TVe2J4JqnFCrSab
BjYBiOPgCm5zDHPTsi+/Z6IcRQEbWaKcB1nLD3a3zT4iHZETBk76oVkKDbdRxsbHr8RPDtLxwZBH
lC8njeOJHaNQfAsN7XQN43irvhBpZJAG7SYqS498YwfZsri9H5jNjwzjWs74wyWe85keyJ7A45Wt
gnTMndDEdiEWFYzSubup2USWW92VS9Qf6vuMOL3SiefYV/EiSaLHubiioR0abLeCunlml60OVpZ7
fnOaeoOWoYHNBJtzx4cktE+88Bxv8GEqo+EjxY3hFAXWoNlQ434w1S3ErzCivLZ6fVo9DHUkzALC
BRwQXmpcBSoEK1GBmqa1btHV52MG7nTvw8RBil42SgyzuMXJEQmpWkC+JXEQV8GwsBOuHQuEroFI
dAt+xUgIpWN3ahPjVCkeZWvqK/vUoWT7+bpNm1Wuei5O5gHfNCP0nX6IWsWBY1lf3qOlgb+FXQVF
49nFbUS/uHGxs4RWmPhbuRorMqpNz8Z7rX0s5Kc6oLbbdtUucC7cTATRclSgHrLPgN1WsEAmA8Qv
rk+cA5CSY84TrkOlYUVUWCMAqKNVRjD2z6McIOxggkbuE1S4gUCq3Y5KptV7kJECSYCUHBIfkv/U
b4e6iGFVHy0gtgBNny7xwPK+ioiTvg1c44KSYPBdRzB9267mWbqndBwW0cHRZqkbJLojhN6GgE4j
2jJCP2+tt/uiz8qYSEzAhda9sMD0GIYAoJRdPgKjFS1KoA9TR7J0e09aknSS71gFMkfp7F8lIUGA
84Fwtud/h4gXJaw1oqNbSGdee2xTxdSYMeIwYyuimFUOH7LX+hXdhy1krKjTLsHRu6pKD0Cv3Na4
zT/PAZpJsfZ/d0V7Aami5O6mzWEyCzb/67HoNEnz408sBZ5y/NaFmJ/SO40nyD+5KE4qqKN6+kV1
GywGPNP4puVYlWGCuLvFbeRub0rcDyPVDCuIn2FCPnmBMbpJy/ypTcF1AhL+/NXqpDoHYTaD0qUr
+n41AXY0dTXUhw4abMfJvbFXWGaUm9ghlG/Trux8TizAmTp4tZqNqUe9sqrd+k3vej9EYbAb08gf
Fs+fgtEsWXGLWJto5puHWaCBL/BSjbjE2WZnNrteuxw5MGooA6LkFVENu/bLFcnnTBZmp87Mmh3H
j3ZoOBqie/5YsOYwNndbGecJEamz2xP6juJQo/RF1uFqMWOoSKxfnBqO1spnrISS0PBPGwV8G19P
EFqb93aqguciVWEie4dWJ6RnGlOi0r5Vq4T8cDJefKvYqHVwUzPAXxiOox7dQ+/EhO5xPEzvL6uy
EfjGcd/Bp/SLgbTTnNZSVz59bwVVJtTMXU717B+W9xgrmVqDrLoCWfpEUF8R62hFCN6LJDoCKi9X
UBcpd8mRPqo2cDgyFdwvf3HBNEXu9XRHHwpocbL5+UAcjOP+CO2SvLahseKU0zmhwudqu2YofW2o
piflWxrQLC7kV62qohLPg83vqpgTX244ubu6TIM79XFGZwf53IY3MzElolNiyNipTBV799+RuIjB
StSKCRpTHwbboULlwsqO18S6HxdC58X0UGE74+L3YgLrCEWfX1fNvrnvHXNgMX/kw3QQh+v7aZxE
gKIMc+AT85NDiI0g+MMyvHVOSqdKPN34TvdFd+kgMt3WlWnW8fA81tIVb2BP+fvVMCGHiMS9hrsE
z54mcAzZ9U74HKWDVvRJ4SQ8QTgqnJ+EbyVlyIqPj66f72jxacQpczAJ92lxd1lA2anRHgzd0MGw
OnmKabWrSRJY2sLMp2vfow15/yS/XFMzpePPsJ6hsm4nEzPxocR4NnU50wmUmmGZRPeTPRcrtAPH
0rHKmuarfdBek51m2T6CplZQHRMg3iO60Ve8xayTlfxNwG4EKGazFkJtROhn20JKhldAiA6uQlOa
a92kuwA/YMlywdJqcIzdZ7QxKYn90RnHxJH/9J612rWKPR3Ud9vucYskdfLYFjcabwZ9OP3fpiKe
xGMnbnGr0ZMwnxvZQSVEFm6VTBGA7qQhsfMbOR1jFIIYy4L3lijTJoqb5UTB2oIVOOf0tgxV1xZc
3eKlLVqYslDMLRm+BexqxUbfSRqkThv37aCRFwbB0Qe5lsczCjcD+pmUWu6G4ldPX+FSh6Vo/a5K
z3xYV2bBCLBLjfDocLQ4mn2C6/biaq6rjgGXwTu2dHkmt85bXoQkvK2bK9UmUneIaoF0Q2S6JmHp
qWD3Md/6qW2SLYpRziw5E323NrnRgAlxxGCy2QlfDZipBjGPC1S8NOH14YVZnLPi2EZIZUzim5bS
mZ1AAJvf4XCAutX+SPGXFyLaoOVNpoQ2EVaPgSVA52iZxqUslxY0WcBJPutcffTDTfQMjnhkIjwL
vabWnBMqni/0V1+/X+Zi08mhrLOHocAE9b/7FdAIdyD5WGFTS4Bdznx882WY18hjm2Mi4Ptf7s/S
eafq1J4OZCshY6cwt6IGRgWrLgb5kHlI2Wfv8CrNHIhskDu+61PQGIFst1RjLnPAKhh99mAZISOV
C3E1mo/myZvo/vf+PyvCAFnHxxHycjcXCxnWwCvkdMHfmHclgyQCa4FAFcZCKRzcTeORlqgIAV7y
p5227xKpo6wh7kIv1lDAUFoL3DR4af9/Cj12J65ifd6QV84PC1w+CPmwrmNTqyLgVaieOPkFuEP+
WkNEdh2DKDI/W4Ln9PHqxUFCdXtLnOI9Fi59iwq3foaDv5du4QM5EBvIt5neSIcmigcxhJ0O8RQg
M5AZ/jElEjkyoniSOTZGKmTX+5NRWooZSYcvVHm4w6Tt3LS+1JukBkQ8DEx3Kxn8mIL/JQV/kGzb
UNjOqvR4rq3VoHQHbCrfWQrnSbI22QYENh+QKCA+TUbOSKPAoJF3MZCP9W4AQwLcF1rbHd37If+2
MLDwdFUSO8frV1MadskBsPpLDVRhEHYt7TN+LJ73r3Hoh4jQ+rk0EJP086tXQPD7v9h9OsnlYUuf
+wsWkmzEkW9Ow1AhaNsnugAiW4suoW4oLJ4aQV95lYLnhxs1tMA+nFBKSk4Zm3NhfFPQ2vDu1Gta
PVawGsAhVuebHIWdRsvh50Vho8lha8tRZcMMZwgKkV7JFpt/gMywYTbzJoIls7NV0RxfC4I6/Wd8
5+mDAvjq8pEf4LPnzL/DiX5yVcR7FyN8hTdCBJEUw0iLCXIafk5U1Aqc38Hxqkb5Ot0t85RObfe2
LOtDIi61q61JqxYChnsc7c+aSQnM+4FuSVA2MDHy+w/pHMyGADllQ+HSuErB8rorJGZHz/TA5Xa3
UebZ6ufWY4c0Xh3RXyIAxF7c2d4T7o5kRkHN+A0bJOpLzyikqbGKQ8Co97g/e3o8HMWcMXhxy5At
dVgPn/c/DENR+qa+4ySIB9JzBN/Tzg+qJ8An/P2X6V64WwlgWS0Hi1dgXrgz6C+oR6d8U6JuUcRw
N/TQ6Kh9bBl/EYfucnHilxkVpNtsxFgLTT7OtnEsj7yfuVAdlNT0+eQC9L+FkXLlSY0rpBPqbO+4
Pnc5rup2YiHOegN2px03HjtMnKyeSOVmV8M3XqMRkIXbSdQJDSftJI96N48f7GTIl9Wtm23sqHoU
d7cm7CPF0Ao8/6kwCSAZpmuS32+MkgHqVod1DLbzUVeD1xw1/sRIJNcRXigfkzq01woE/5AzGbWK
IePFK/eVIj0j5sB2lGbmym6NOOL6VlwmUhg2gxuuQLMFnLml5z45docjdRSLg/KuVwACvHzbzK9i
mWn1b+LlZ1lO7yXPXRHw6witqaxwmK9jTEv9qTCnJs7MMr3F5Jf+9DTbuS6LEdZy9Dng35GEHD3s
vmM/T2zQYPIl27fxKq7iFil9k0rvxCvdg4YViDQ2tmiNS+nKyFsMJxnEQJA9XYNxRhjIz2IT4rhB
RZke3nJR+Bxo8j0m8xGVDkoEIoD669dJSfL9f9eyN72oYKt7bxS1sNeW7oHSqVI1HaOwfNBgnJcr
L9xUTjqW8M5WYJaDiHyb5bS0rKEf7Nao1WX8lkjgsT8srXPw9cPZ2ZYkwYYMPaWfFspHE2mHdr6y
aBhft8dLOjCVvhKKxwAUImOtwmT/4RkIrDyNO6kNRXtIZrI7CwNloXvd6KwoJrrdc27TgJnzTJB5
u38nPGxkEm1XpXJxrp6PWhlXcFBH8cXVnoN/z2jSCoXCC5Ob98ar8TF0Zp9iEvSJa3j7Fp9JEDXe
gkWIrSTD/3YtBairfnV/jn+OhgG2cDrGLUaY7DhFJBytoWVJjJ83AwRudkbD0uP6SEcsvn9qCk03
qnfq7CvqNCVr352aIAxtFtLa4ZjscXBDN2PxtX00oT0tQ579J6V9BHEWI+la2KhVtOouZC5aXcip
HwFwvOXkrwpN2bIx/c7idnEOVXVn9Vp/3w4HGwghOrxRHaPXJmPAI/JB4FTFdkejfZ5IqWF5z7aA
galp4JszcTC5tcmWFj4J/i/Tr1OhUxX1zJ6A6gKXjPnc0PHhQbHrrlVDmD1Ixuuix9/IqK9dsdYz
wNOiOMhTK0u28bBe8olx8/pmi9b9Tiw5JuSw9/+0rMLttjKD1PHPLrNBMD6VXZ42BbiOUtXRXyeW
zmeLKlc+lfElb/KlX19GqdFJg3U8KuB/XeLkhlloKuPmX03IiIX8gOK+MlY+/zub0NfF0j1ROEQ7
ydnzDAH7cbBFMXJp8ZZcFWHgRWou8C7BqSU0PPUwtWc+dHT3ggpo3v/bP+GJk4JW31CjGVEn6rIO
HigS7q5rLy5tHt4L3tLAXrXeeHD+CRf9CBFzDdBKgrL0xUhSI0sn9zmfkhalBQUl2wbHYr3eK35k
Dxtjt53PMa4Jhrg+ySDSv3kLcLOtyOzQIQr54GYnarIac9Cb+a7hCa8eRMVyQI2hd6gOCvAbc7Dj
qAl0GcOsArKXEfwJdQZdaycDfomOC/TIBCIJHHJUjfrSn4Z/nE3gUR8DCwOk4MXpWHl2TdFkUdbg
IAKLhzSPnWbIFYXO2uFYdN5w4+EB0CXlPBoiLDvC734zPUSIZhFGCSftyaowAP5SrWiAXDjwWfbq
IZZPgemE6tdfh0P6yepIhHMJTENW2Vy8P8mtg701NQhsKh8F1+M5DhmJDY8sd943RZuQTJnz3b0R
YokXB5TEStq9ILt+A1nS4dmyucdXmbZRr2aGtXhpW7kEnqk2Rlbgg+MNypu8xw0fTUYzPEkX+/ux
CiugucWhX46QTX9oNm9W0qMz8vztMoFIBVUyo6H+lqrzIM5AsuZTD5ubnn0QS/7Omq0vI5u5hvmU
6TUlqtdoFLTf390qbEGlzdEi34c7ROyUPtUAI43Zijf4btpQRoa3VlyOHTmlAV414H7HGmfar6vA
eI7cJxNLPpjHPYBzLDVB1cyAtguOLh7aW+REOpcGMfF5x5Vpr4xLwQmlT4LlIhIcwRA2Zu7XeleU
Hhhmbq7TCQq2IaHattdJ72YEZrJGxVh9uGTZ/B3ST6WLL36PQsc36YjjKgYbU+Ew4PYdhaNKCwX9
ZuuJySQXuo00dvTHaXwL+ObQMA2xJ8jWTh45Ys3iMJQHRzd0B6KMzz0nMJjoV49aW1ok250ijLnT
L+f9NoZAs22nbyK6mfpc7cC9lfL42OQS4hoWKlk9HjqZz2SssLrcyLPWJe9hYYXMFy3ZmksD0aWQ
2VSP/uFPx7G9uFPm4TddQzIZNwD6LrHzqnZ8RiBieKfZCZDgvUuLyQQ8l/s1cq8rbH2wznFL/JCY
CEMky2xn+8ZhXAbUSs+x7ntv9ASxYcpQs8F8xq5VpGCPjB3UPSYzZEvcK9YKJuHlHeSsoxEXHT6Q
1lvEYtc2uagMHckWjA5BsOc6hLrul/AJLcCdjqAqzR+sd4h7sXnozJEYpP2HdMnzZCaLsHL1huBu
5S9y2unLlFx5cKbyf41fCTYcMJ6Mgv00ke6QNqi5q46rAn+I+BpRoJIw6zIxuyNTEWXYjG+r/rdd
8/4ASMy7CrGz2iGK4+w6HUJO/HXTTnZ8oD9oaN4Ni8E7js8yo+NVYvZNO4dy6R2HFjjhHGlFhKrm
2LXGvdkH+ftL6RQyM/8akXV2XTY1tFCC6hJchoNqACkQl+NTuesGA025D8CFmJw3m85CR5qP+bw/
/womeW0F5MeauyLItxYgN6AZmtOCihTtALP63KEUU6ZUV0+5tOhDm4128nSH+CTMOm2z/PcZ06vA
q08MMLbkCZ3yisYgxWcvWg5OWgDbSNirMiJ3E+uBqM1gj3314mx/LeDGY/IT33cP9oNZ2CsZ1dcf
Ber7vSTVA3qwK3rqInuEvH1QLO8hYJgIV4s3lii+BTmBtC/1ZOUkhibPVbMY6403Vnyn0J/U3oLA
XkiR2b7ERt1fHHJvTJF7sv1n20crzM7CAk10O3a5ktFYjRS8yh+oNq8YSMgHM/j1rRkQ3O0kUikZ
a8LFHFTDhY99VEwCBL7Sy5L3YjtRCIltaPOs+CxDAjjK/0FjjgfvPnc2RBoCOKbDGCUXs0tde4EY
UA57Rsza5GqGn2lbmmXmw0//XLfRuG+kxQBIHxadUbjjARAlsuD1o2d5UpcxxM6eW8iWvY6TLA7L
8NARNWu8wp8BEiheY/uAnugeQ5tUWzjzNQtfJV3Adplz3x+bqqQLCvXT5cLu16TOQrvsKEOVlD2y
tFJhN4jSQ16RFvOYxqraND+evAhLSlDNj4977FAJOTgeNFrJyluG33E5aPHNyYoyquNEj65Cp+vF
inlJUH+LjCRnMfaNpaEXcyAdhW+FI763+qWxJi3Leii/elpAkdlxKzWlAiGOmW+SaFKByni1CH8U
TupJd8tki6GF9oswJmYYhgzQdoR9RCJ9v4ROxeAOXHA4zdNcKZxcPzoC2mV997JS7S/a1neBeDNs
YD2r1fbKlRjdAYO+J2Vt1DjVsLvh3prjIbYeyxi89ApVpgzY317VYUO3sAC2a8qp5l0l8LOdixEz
lE1SmNd5Ddl5kX14sIEhCwLf79ok6ZmtF1WF3/18ie3Ql+Kix7sT1UrGn5ti63Yz4IuOPzNIhx5b
hREQW99P9zLgOAf6sGy9iUMq9xE3VJXPvRo1z2FU4sZ53/dAqMCUChw5RXhyqH3Gj9tW16/DTSUI
o4wXs+EgvtPs/CD7kCXIwAjoV3LlmdXaBv866X7DrOYp8nhOPfhGcx9mcm1PtUerNB8/LFSI6me2
VNgcroL/vaiT5OQwulcNqVBxm9WgqndBvGp59eADLYOPqI5Qk+HAOXusubr8KKN31SP4P+n2DVVx
f/MMmvdpyvNn7//SiGuopjBIDtk1AVLcxzEIp/qEWQaoRn/y8LzfymgqvPSpI+/UUtprI35Oj5R2
tGFLvINZM5X0Deo/0E7bT6/VLQGyBUIOcOOojX3VO149kQtU9n9NxJRTFG11GnHY/28IlU7Z42qQ
TtOXWPo/nBbkbxA/3kYpjpELMlhTZlMkHNfpTadkpbIVXBeUGXWVERZB4nkXZYTTgJfbZk8xRIaF
x2UF1Q1lw7sK7To2Fif7N43489yWWgl3QuM5BV6B6D30Mne/LXE/voi6vd6AvLOCS1NeO2KUtuCs
mXbjH56dKLTCJtmwMs3/PLJ7YE8/U7VpeOmeokyJpRo2pIlH1dQJ7k7pvB+elFRg1yX4YOMhdGBv
RpO7ebQielUjz1oV3xMvPRx3vxSToJeEM0AkDur29dei63Y+X2Y4E9FvtoWPWC0zsAv1034ZZa9b
kXeepylV7rHSw/k72jmm6u+SG0heu2BpJvDcD+EH4C96OCA/p4buNGzwVsPsqJAU53vB14UuNP1M
TeqfendS5vrene/kBymVldMLU9P3UX1Fk9GAHzJWnLQrXkZhXGG+o4ep6K8zPp3i1X0jxztk4D0F
fiPNmnPr53Gz0RN8ePxxHqRzPspBW5bmzrHiKtNPQolQrtmlyqRZ9h2IcwVmEFZZdd85BiED55A3
G1tXDto02uhxMXEup/nzFQ49ehrSCsYvhEXnVSvd7EpN8AzyIbg0IS0EzeuwtW1L8dzTuq0iodGk
ustpKasYheXkSaCj3Z6ycgnri8VCOEDp/v6HWguseCz6oXtzUE/VjNpuUpsVZugDXvLxdczm7NXI
DsAVl8oCxW/MEC8Qn2Sc3cB+v+LHPUoT/4mKKUFLLAP59M1WPF/ZYvjtxzkwLoGY+Rjwq2n23k11
oKyQrqjvdKDMpvr1EZ+C7L4vMxlBhBqXvckdDRs3SGCTLCrCBnbCJaASm2qZ35w9aRldQey4LIZx
nPzG9hlBzcr/VhXS6vCyk6qsmZ44LNvO3KGCS5eOc9A6pI2PhwvUjIna80J7UtdRR906PPc1+l4n
peiYk2QkP1znvsfJvZGrHkjvpBYTgR/OwcRPsMmP9maRw2+gVyAieCDIe6IeJR+JUrc3NRvha1Ix
1r+ce0C9WFhkSBkjq9S5DCQHgZCDa9p/tVYtbmCSI7ANrYW362VfiKaFw8pmyX4HoxCEtz/i9vbC
s3ARdoNpITbGQ6lCFAzoVRXBw1xDcE4nXzrPQOIiDsARnEx0BGGT+TGG+5dSbOXK24VT+tHBX3aO
t1ZdDF+NbHUekluIBrxwhRtYs54y29PfYgoaahdN+xwmH/O/fZa4cX2BaZfgMDDrv2h03C/Q8P9M
0hy8nMlroGK2mZM1xmxNqAbH/HJD3nyAUrPT6AVSUYaYURBLPDN5A3rixU5ikDG5COiof4/FUNS8
grWjy7Ymv8OOxw+MywR8yeRVy+5aVZ7aGN9Vjutbds5M+4wxpzOXWLJp+4Q84SmQgFGSOptd7J9E
dWAptAalG7TxCmLeK5HO9Rp/8qBh73g2FJDG6jzXvWs21M6rokihI1DEwSn8z8kFkq7J/FJvzgaE
s2oniO1gC2al9ri2k87z6+UxWWKJ/LyBEkjWaYq5emkFxaSU0zmJJ3bPobomfbTQ4V8CEEnLcXfv
XswNdQN4neq937FUowS2N8PaMnJjxBS/zGZX+69+SL4TvZBzmEcOpMYXZ9h+pvKQl/1H+7JKyJG9
jrfei2Ma5R1E5BiKO6Kl3OVyUTWEK31zjiEvlJ9PZl0U3oicRqKwerlBRr5syzHYxDJqQTCrEV1v
rEV71d1zlvHz+RPtvjmdG9FtcCwnHW9Nqtp0xuge3EbzH6j44w7cqp7CKLPOv2V46ZACdsnwSGMX
1+wBXyGVSMRe4GFKzIC1ft7LfKeXu8CNMOVyDasPUJBI0KmfIDK7qqaer1JT2XivfIehtL1Wou7P
KLxK+tKv8NOpkZrqawxBKSxfVupIEq2P/AnKVzSeN/9Sf3WjtR5/mc/X+ucia/ejdZBlofsPWekr
y1GcPkpMKfQIr7HgUXM1+u6G/JJ2q48m1Fa1NGPZZRCFAFUDRwqC2N8KPTUqsITS2yFQhukciDWf
FxCXrN1w+JjVJb/SJFEQA0wSR5Mm3SUSwkjs7XYamr2ubIHJxjZwcm7F1BTgCNXoFNQ0eFnDULcm
c6VYa3NzrQgyrcBU/CNJcV3+vjXK4CJ0GUbNIzB34uwpGN1Ie7e4gArPT9TUqhWAA8LK+gU2sjXf
bxfuF1mZK206YJ8Phi3MR0LOuSo8IFDH7ru2CfbkLyPtU6alq1/3qtJlXKgrYZ9Rq+Z1NMJuQsMk
R4+dWBHpj5JGCr1+8b+ZUc1YKFQtoycyob+NqJjVY51fLND/bNwzfc0tbZaxqRVunPvom+bzC5dp
vICIPB7tX8z4nhIKQGZPUB8naadeNHzykmkdt+Um0F/jJbzLGnBZb6KdAlrmYr2Ycw4uNYuM3dKq
PWQjP+q6qJcfGDMpxcNVKOi90bpQhfGEb36k2JOra8JyJCuGXqIEJ7GJRTM9LYKx6WhF6ZHbKEw6
yaQoM1VK638EwYem+jFFsFGPJgr2XHIyyyp05GaK7p1f8GPeP77ipTA3l8yr7XOnKXh8UmYjqX5V
LRCaDuKRbAB5w71/nnWRC38yXfa8MiXQKrKBBIvE9wqPs/EK/YY0LKjQkBrM7VThOTBm21HgLi5R
ot65NZ5/dXoRVHkwDYvg7zo/M4SyzNUZihrNbs+nASTpC/zKTdcJ0BjArXNZ6E0N+sFqQXYF0oiB
CzQZ+cMxRNIuU1IcQudoPxyfP0bsA1aSoQ91d5ZWKsK5SlLULS/AYcIB6ldPNJtkq9HmsK2b3PLv
kz+Wjfp+wFu0wnCbes/yBfcSLnwt8beh3LUpW2aBRlw0cYlvtle6SyVm/QvfuYECVhMFyGKfBSKx
nvJ+J3CpEeVFwQx20BUidkVCgVXFRp7SDaVVBh33fwnfH+CL5Jkc7NtqQLovNmNbJy6x8z+jQ3yw
q1O66x1UVeplepSrymxxMTs0AcL89H1dyGPO+Y69UONKXuengrwohT88SNld8/uKBseQFnFD/UB5
kiUBiw3pYCcrEVmx4NsASNmvW5pgQ7Q6XkSapNoQh87cdZAL1mkBX+KIEJ1sRreW46+SGf5CzZ8A
/OOKuRBOaTJXYtcTlFW8foNZXmUWl3DqQAovrpyoKkkpgfZt39LI19LgCuiIEBDN+NChxrqnOTbK
3uHyPnwvec+Cjq7zKvf0aYyfowj3h4x1WY7iPoD2yBPLPjKMeMRCLthKZH6qv4/rlgk78X8pq8JQ
ySLpBLRuj9XrV6C6TdpQR5ZW7Ns03aUmJcjUY3cCbhPJ5BPnfk86Rwm/z6nzDj/mOKr2r/a7TyZC
QOjyk2mce4PTmgsGpQpqNufmUZvjkXLoHF8uQjFPLyfuheDZNXwelvSpCJnZTyUtQGJgKnzpHyQO
XiYdVWtRLbPxXGnfmIAlZQqF6ubRt4v24MlPf2EMVlOOjs9N362dWV0SgIqXzzdn793Evyf++9Q5
mo3L+kbb1d1aSgJknA/7UZGBieKLJRsS6ZXZpmgQHa09yfDzYHDpv1f7eG5f9tB/Qr5wVUFRf/aQ
GzkF0Er9+nILBPwh9Mor17Mj5PgC47cwB7eX31EOlByC2A8W9s0I8b3z6fyN5NE8KnC2W5JFxMwE
Whh7uWUauznv8YA9V3L6rMvXpavZXvSfnNzSVI9eBWpTUmJSB7FHFz7ZMmXnOge+TA8zaVWHdpzi
QJkMhBAHpDDV+28kY05OMZH7qTfYmH0ALOb+o+DuvEt4mX4sMPaCwFzcmgNYBik3583TKAlOgu2m
Q4yjNvfiebZg/zj7vhQVKX6X3j1SRebDVeRGK741SPcuGAV/HcdEqDsn0Hpcigi1LVm6xUNqXlXI
jKHgETEpxq1ZZpbGl3ZPzxoO4AzHjr0GeAyc5K2FM8ak1cJzt+lbZWmeYSHLIA1mSUTsXK+Eqfhs
9mcZWe0YrRcVspGisBCFRow7eGibhiFXcsT1jx9MvYvtTHvFgqMiiimfRI6kprq5JonRraINKrZp
VI84zi8OmvVoTRCiphyabKHGd5T9NucGtDByt+Sv27aipk5OtPpqBZyuhcYTyZPYxwvPJ9AH/VrK
OF8WcSmKJQbL4Xsi06qqv3IWvHjxGj7gdVvRAffszpHufg3hOJc84zjpzde3a6iY11eZo9snbpFP
JaWkaT7lfDStACwx1EwRsNja1n2EIQaJ/yCzWsZLtHgkDk6StiUfHazxYvQsCXvLWapBO/G91lfa
brSxsgdSYeDSwbh2MsrheV6C6rYNmv3uefeowMck3F4S4ngoGoh9Nl9635e2uCTtpfaNfzNjYjw7
C0w5hGSV8KMbk1gNydpNo0oJGWhBn3Krolsr5WP978odPFdC9qaTVvHNJhKJGiw7z1Kz/z9pvFHo
I5hMdlTqbAwlGYENRLmBqzo6WZJxJXUgX+milaI9y+kh7DIMBTXOVrQc8M+1uafpebKXA7geXR0C
wl2U5zhBizjpnITt+f8fI+Mc4z/JxlttYB0aXPDjRTn4dDfO9heeE9c1SWlAwdWDOYwtkXhI8GrW
eVGAfnf855ZS4NhCBoWH2sQl0Vx9LskMyletAEPdBYbRsyAxBzh5sT3cFMPHmEmC8cq5uT8eJT1i
jgstHfWCNhJPpPGUmShYCLat8ESdVTfrx9f4B1ZKmYvGpJ2tRtHP0ZGjLkcfJUDSCRGTtx9Asm91
l8PbCu1gzVDOzl3KqJ0MremtgdfNqCghakXtV/Qpm7OsGHC1A61KryprDVB0TSL3ElcakDDsvnGQ
T/LVPt3sX8bBs0T+RPECjH7q0coFcbVgdNs0WDwkh8RIF6vVKJlTRb9OPmmFggvojt3u7dE41PKQ
aklwnrxsVdSrPMgHRRNOp0NItBVw1id/Ane3LEIfNoeDSbaYz2JtKDzXARcTmoKgTLpXGyYB9kt8
ns6PAndXN+K0aEPLGbqhNpmFpQeko/NdkBIF2f1BTf+c/BzK/+fAHc1MDcnd3fpOtcKbOmSZsw6x
6f2gU2CM7QS/qfuTheVCjMaXGp8sSkS+Aj4LDQKqEVxYmpFZag5few8ZkUVSO0mCr6zaI73UjNKa
WEVOgIE4EgCXqgBb3XSmR+PqMxsFSfZmPhTs+ndbPubE1drHrhx/NDhaDAxI7889aVSJtlxF46Tz
KY+/e9V/rx8rcRhpD7O1L+Qi692HomzROhaYIS6V+POPKuLgyL0iPEbEOeMauCO62ELKqdhbuZK/
xoj7UVlJrBwPG++TfPalDVv663xxKp127Sz8nNatGA6scCUM4Spjjxp7oHU4Ibnb9EDUX+P0KoRA
XtPnX+rQ6LUGWNUqSTt67yuAwuvWtsjDeEYWHV6VJvzZ1CBqpb+AjEyz6f845vsEuzNcCoptiet2
06dCyaFcNV+J6U33GTBybhY4fPjqVek2dMi2weAM0MlkAZ7itgYmSxo/RNwTvGxVkNjpv4sXn5/5
22wLbIAeQWJKNoJty4BdICqwGAPjftpFBXTuqLnXfan36uOcb9xIOBhgXevtBh3rOrcuPLcQhm15
mp7j8WNVKCwmy1UeqvVr+SQkdMlD+ibxby06PceoOzeZS1pN9SGkRwVWaAzSkHUtd6F+fXoQ09gV
Njj9VPG5S6YtQ6FaCUuW5Deb7XN1/LuC63I4ZY9OIFmVHbHjh6hgNXpez2zANV8mp5rMA0A6xEYH
dIV3bCMublVT03vaMjsAHXM8Q6aHcalpNy/VHg5UcLEDluUTUAjUK1oa/hRl2YT+ikS8SqvaXodG
9XV/mk1W6xu4msT9UY5cm2x15H4otQk4z26m0N+I0JmreexQEY7VuKfsONifbDIOLCk08UW1JaGL
aYF01aVGTAPZGzQBzN0Bx3cl6UeSuVC1VY+hP3ov2Dso2MXosHnZxz7LpjmBJDR82N5tbcY6gehx
SJrk7D6GqgnJ1rOh33oxk4RNA9kdFYiKzqmFf+KmU0wW42E3kBQD6rjp7iFvdqa0qxawuPC6x7eg
ICWKY2XYU7AEG/v+uEspojIlufTu6f98JPQE4KPlXxmB4ic4nmmX2OtMZLijD0UaqN49xgsdL/8R
bDvd0mbwxUzKm6Mp2W2S2j5A68i6cCM4ZBKqbMYS3WKnnoUdypkDXycxo2bMdFfkra3d0gzuG7i/
YPIJTpD38LDpnsTLBxpoxB1gGEMB/f1CFq7joyLlUfivl+FiLT1mbbaBJbsVsL3rfidex5MJjvzy
XyHVsUKdmApTXDecOkIYzYb0ZP7t076Ji79HDsgcDPkMDNLGYvqpXxo3sVA4LHnB3/8DrG8ZcQn/
cW8pVd4HQfbMhffPu8GbxWD2NNTisaevE62e+5w5Klpls9xZ703SCKDdv7I2ubYuGf8LGgZhr38T
P8E+Rbm01ihPArC+hl5OzsZOSCz9lTQpBQUfq4WK0we8oUIYY4UJ3OpHy3eaRN0JdRtYV781KSTP
7/ihtzw4xfY8KPzry+Nyb5zhnW/jSfQc0CF+rl+yH3Sik54cf1I3dnPWCzzJ40r4yAfdsxi6PkLK
QZM87aHtdjZEv1GEhYDGCuM/4NlCaw9GXhybArqZobD7AQbrPSFOAEA6FqpAnw8RLDjdv3/kG2kd
+4ThtpuagnByyCB8JsZ6P0HP0vUJy4RtMODhXV3vLmtIlKoq0d4wIOaAmd/EZCr/7mldGEMXymnN
LXG5DKspLH9gg3mmevG7c311EezyAMbaQaDWdYH1YlX3pROxpvfl0qTDfkqf+LbA2Opg32X2m9OQ
wd+ez9amUxS7+1eIuEkD4z0wJnY3u6dFbvvnn2bayRtOhMOXULJqG6TnDh8EXd6gTrSCX4hEeWFX
GimpSDqvl8NytyahkF2PpkSZfynBOYiBzcXkpe6tjeJxodPPk6ij9tn/CUX7wvuhzRvmgeFlvYTr
ExxZruiOQIO8oyyp0nrjz5yFon5oU5/gaqNrxc4ZRh3hftATvbA1GOBPSXYZMTZWpq8DSbpfGnQF
eAsXf2Z0bG5LmuXxCerHmMgWAreIgLn+wixCr2DeMB8RU3ak79ssdztzmDk05FVxmccO6gyOXofr
/3M2FOJmAEaFMTSOJvwdicqHBD2mJAGe180Qx9GJT1TWFNew6yyQIa1MwGEgiCeFtq8AT/+vyKd4
emO7VpCY3AhlCU64s3UUL1PH2DrH/pE0ZkNJAx3J2Hf5edwgm6IdjqVyTuWAqvBdRtzkRVMLM0Fa
t9GV8nS33lxZQsNQOjIVSbUvFhSvoLxkwGhh4PMSRmzi8wjHr2rcYF8ohKhIT5AGLzbouoh708BX
1PgXut2OcWY2X6vMMp9L0unR0eEkKtO98noAzLO7djKHNKgmpXKXFwtyjCL5E7nlxw1Q+aRWNmfN
7AAqO+Uu0Hufqo3SXPfi1Zs4a1a63Fjkpw1iIcYQxxuh0itqHM4mWX1du2yWNCv4rUabrewP0UAh
dO8j1lZatIviv2gkagtFpdz7M+qOK15rTM1h5sRvbPdhlNN73srJgGpsM9byJrXuaEKiWUaUQpm8
TdOPYQoKJgTU+WJkfeWeTD6qYh0VQBfwIjfaiOQL3fb3p1osaWVqTlZCR/EhqmrVM2OlByTUH/aK
mKpVnAN4GrRHsuBeruhBpIrl4Jz5gGicvjoQ2xfYKYvmuP7mpqtvkjCYlizdFOxiAddG/9GENSFX
YTFC48zbNHpaRjzY1ukST3dQ01cTokCMdvutURjBbWY1UL9BJkxv6JbhMuynqVqdQI0xdN0uNbbB
zNlMBw9jGlBG5LQeuMiyH/vCiskvlhoaeA/EbonSDgiIsoiMsxaccfAD/83z1HHwTCvLojhzpJrz
0XM0Y1A/ZbTrkKRvKtgHJZsdculbqsR6Hwy//uWwagV64iqHqDtrHn40qetq9ZsK6LeyCTVD0L0n
txayy5IYty862irkKyJmYTkj7Y3aQiUJO0/5lvCvS6qakv8LADLfDexT/Wx9kdY+Hy7jyBJsNCks
pjHVKMftgkXYX7OL7xc4Xh+L2Gg7MmHiFO9wnIKjcl0WHjI9stcgV+k4FzwB+k7xKRYoBEVUXD9W
+28g6dOIqf7VvY0En4o8JBGkgLyBXxOAG9UlFPhVNhs3CsHjDf+JXpTbAi50QRtP56W499KszObO
3DtrvlXlORYNKdGY1U0dEvpCffPj1e9QSOd6sNbhAax6ZVf9ecFDyfA77W2Eehz9WUfLtljOUMGF
PrxgxnVO0B08SWSkzU+UNpiUOrPodD+OYCZ43G4d53PXi7tFbUROCM66Flm0sBMSkFd1NDutu2Ny
mcy5IiIV8eFIxgnEO+SDNEAUEjlyB42Df3ytL5wcscRZukrIxNMaNTrvqoeirHjKZqO0u4p9/5H3
p6JHlsNii1gx2XzNB95LfaEzZ9xlJDqLoPaED/EmOEH1cxWbvYGN/mz1K3TlVJKeCYDWgBpYWx0r
EgkFa9oJSvkVgrhPZj9ZHerDP9iQldVMZIBzDePGBGM6R/DVegXZyLa8B0hQuVsk07x8taUj7oCO
34CeMpkLjMB9QcOWB5TkHGCxZUMzQyXLnKOH6JINlG8eBRoV4TP5jgfX9mV+6ecT8d3CPO4X2xzR
DspqzmI30TaNs388iJJBlihgwOy5uEO+5f4zrETY3aNp47MOE7wEuA+ZsevqoFsziBYIs13MasnQ
63K4xf+InbcqJpj0wuafuV0NLiJW+CkdJp0qhVcuy1CqD3KBNV8GmZ6c0u4BqdoRLckjkuMO0I+3
8gUH5h0Z9YZzPo18uADep/4i96tpAl6r6F9deWdvnvAlYlKlJIAFPkzm63Hyv/2BURI+HjH7BFCU
D0M0N2Hbm3SdYLHaG7gg1tSgjSACWWm2OdFcJrzMrL+IMlEprye4aPcIQwaCZ/Qxzc+Ucbysoe/g
YWQmXmu1rRfJb/sjf2dbY03MXHzPgc7usz6i1kBC1d8o4z6Zx5L3+ttLGbZKPiv60CL4CSQPScII
+HFyvM2yJ5Nxi3DPdrEZgvWVFSd+J63RdpNq3EkPmgPW+VwyTcsHNrWH44bpbeBso6rK4drbZ0Jn
exqOo7eQzvft6wR7HYI6UFtxFnvitYjTniEw78kdRkyI/qvzhQVh5I/O3ETsjz+DLjLNzwEdrb7l
2iYeXUle24Szt+Z/sw6wGfDZuY/U9Ec8HL9X15ZGDlUDVTZeuCry8HFNgARwvRfcMNVie6saJ0Nw
vyJ1w1ZmeNLOKLuKkyntLHV2dMVIPkKR8Esx/9Q8P3zPlx0ChYLmu/EOx7jzygwqHC/grjnbjYeQ
+oXM84TBBA87UnA7rjIRA9HrPhd3H5iaAQmQqNK4h5/olHqwVpk5pTrpu1WidDPfuQTTFEZbLr6V
Pb7O9fRx1CvNNtupec9ZqkahjEMD3/5LbwG/3AqM/15KY2jsxzh6sDf+NeFcr4pT2dA9RAfj2kQj
PPU/ZInVQC4bsHvK3y6wQI8FFZVodDXSkU9BTqBpCoDN7ERRApSr3BYuZzm1bwHAwSiB9VPGPxxC
xTD/ro7Lkv+BQbKdv5+/V0hM2/ksurtPM20/ah1EG2Ke2JLo8R4Kzce7MGhA19YCbbtgabrOGf0Q
MlTPZ1c7Q+4Zx3HYRm+jSVBYr4a7h23YPFD+cRdbHPw2pXC+jC7k03Tw8sXPF4Wvt3+qpygXDo3j
YUche4coJua7HjsFKsMSv7qC4sGJgks0IE65HBuXVzoBu4dewGmkgmczaAzjxrMrblTy+vWfkJwj
wQfJ9L1QjwxADczEKrFR+ks+PRRAc9gVSpel28YjZzbY5P8zdpYHYSXYnR8slyOrvIZGtCLLJFcT
Pfzy+B091nWSGhErSzLe9qYNzdK3W9T697XbR4O519CgSGw1iRa90oOgRYwdsU6R1nnUCWjj/U2P
0T7Inb8SbhGNdED9EL6S1X8LfEF1Pa728mziDV9YdZelaxSLkhvFZi42MNuQamcS8jQehciYYZWk
LEXyLC40TJcuO+UQQvQaE0CIGWoqBT1RGOGof69jofn+R4rh6yzJsaC7wnAfRJo4z7MjlmjY09Lw
/a0HqR0qJ3NhUWB+GulHSmYsj1Sl2oBloFuwWuawqIqIm2N+dRDLTsq076Mi274fZmL57TGX+p+W
GELqWDTwU0mtYJ/tuzDNXXJfmgytfAk7C88/Fv0RLzaaAjA9e9gxzoNvhn2mwOVqDzvEHlsTLSQE
UM9ULAG8Bz3w64vvtQuUPkaiEHmxNDnPnPhC8prRQ2bB1n2wgGAVXuHtd9Z008+AbxTYJDZSR9Aq
1lfEcSidI/a3JBiGlhLJTzniKPd9uipEFSTC1Kch93guNY2koJr6fyJw5eDO+oOiiWx4F5po+srk
dKaEOz7nSbhpsbqqJsTxGkGa1uRtqG3idvV4jz2/UYjndmz1FBi7kVsLcojr73DHWbdweX2PQa7S
jwHwxfjtsghHu0pOzBKLk6490Ipu4OXmizVTcHQEq+MDVzOf5tS/bt7BGeMVA6k1j3YKYfp27gF0
cBvqoBA4l3+sTBbIaIs67VDP90kP/XWZ+XsGIOtTU7NJpvIBFz2aqckrCy7C1mdmUIcXND6ap39i
2uYP8eNVK1w4Be2LSltVItWi9fweUIm0nIL69su+4NVzU3E1xeJR4N46br7BXhXUFA1vwXkgFmgc
RrIoCAqNNC5KblpmnNzwQpuqMVqkMyQPO3vUuFG8VhaMXn2p5N+do7PAfLbh5nQRQJch2zOWh/xF
c0ymX/zqO44LmBkXpFlvs1jdGswyLGzGCCsGUONwfBYlUZTxrwmhgY0FFjNg9hst3FgqruSr3bgJ
VUyLSZ+AucpHM0PVHcoGcjndtKfVJl/4dN82tIg5aoq25PubDxxYPuS4U9Boqe9F0ZVnfbt5tBGh
4DnEXqi5t5teAbsRKjpbdxMVgA5HeYmKoeBsPaYg0vlM7O9w246YZ8e3Q3bA0cnLMVM1JXg7Z5WO
65C9QwrpR6IThD7RHAOlLML9M8ilDNPsYG32DiZdWCJ4IoGswSpBbHx9pBF1l+Nz1ESheIFVd3p5
nElhZRfEqVxo1Ml2aRcRvSvKRr0CRH3+XSSWoGIJTM86x+3LJtbW1GIYG6EzKT4WRKET0UhWZa6u
SRLxGLaVr9gucJze4YNko4PtoIXPWFz2OyeoMUImHL6VTct3QVJu+1yPW31TAWGXpXO1x4HB62tC
Gh0y8S51tp76zYXIq74Mb0PZsrY50ulHqbvERXMYAFFSdmZ2tnmyFqwFKHvBMowB6MDgX287ltD1
AG2nUCDfKKqWBhIZ/wAFPwYkrBPLnMm3Sb9RckVeMhyT1laE2VxBnQKpF2uYw78xIfJutCZ/C7Ts
ocjeuP59+hx/kHxPhDDCw/+oNlTNqc7VWEpcNtV+9mIqk0kV+JEPNVeM6cfFmor9npcgbMe3e+r5
Sdjf6X+WPCQ5jr1OxsPZ1WYO3z36HdNNevATt+YH1lJPTSrUS8bCWFb0Wsa8u4KFN21NdmGDH0hZ
WNP/KL7a1YfBwIcu11Nv86uQ6dEkgl8fQBcJJbLflxD37vh6plpfG3xmVQyRmFiIg8qIRFbPzW5M
x/h0huf1/TZ1K/NW4XNjZuKWOHVKWZngIcXIAGpR7rPBxX8+wOoLnlzz7lPYNo/DC7oo/xS5QQr9
jIdWDgzlbZza8x3XNl3uKe2L78ZuIdoLgSiFJZL0C0pu2g2/3hOcgus/ie3NGxBNvyh/f+EyqLDi
WlM3bH3p8VTOVDp0SoRsDEqa3K2zzkAQff/MJRxbAx0NpnD+wkoWLeIMmeEszjemMDne+wU1pbtS
tI6wganNtPJy4ptjUUiEdmgK2So1YrNqnFhNqIr3qjWpNAahXn6LanNDGdOcVrpHrtyotkyeVoGV
R9dXmKBxSBD9ga1uNGrwd9CeMgNkq3UKm3zUGwCJtyoDGPmI+duBIff7D2dwxJla7pOrMtsyc76D
/33gyNm7G5QGm9dFDQdvqcUya/DipmthCExKUyPQHFNJJVTl97jzb84ei4zo25F3TpLA+21FanN4
xF8OyEFevBsQpYfFr3JxZZ3Yv6/PHA9sRas98TEFXx9RU+NMeBNYASXWt/wqI24CPcixtkZcXoac
N1jbbNAx6GYYnkeiDDiMVfLM7R25oOhdp9MrN58mmmit/jWP88UszZbnd9i2PuRmM4J9D1Vwmw6f
aI1AzObYkSHcce2V0LvUB5rCQSgr5AV/hZ8bHZgIyniL3tqttl78wR+j5ypl3/VAiH7YR80YAStn
s5MmMfsoGj6XgtZR/rUKt15lKj+aZ9f3gIqExmdCH13ZWslnuCIgkSKikW8DzwoGYfuYDGySJ6Rw
J8VbGlMM+09fUuKNUHbjOvC4Ufn/db/u+iRjpmTEuGEAys3j78wVBg7XRRc3GlQYK/KepC2tUSaW
cQAwRqRPqHZaOXTzK/xpKkSknUBX1COcqff4XM4Z3ZjJiC2ga5MY+KSbGMdr7xvcg1VGKuQm6H+i
EKEABZg1XD+1s4cTWa0Xf+zCnlcBzPZXApP118iN5nFNMiI/Z/1RLYxEjyQFikUpEkawC40vSle9
m5koT5zO8VaJIlTgE4AgRvwuLcutoALCOFaUtl901YjrT0CVsugpmaJqG4pj36bvDDcCmlMDnJDd
7rfeXtuS4KaZ0s5c4eDw+KM1GVQ2YRdy8LggbnC7Min7kV1LrMKZeSLJc9KmkGQrkD+eJti+5nPx
hrqyni20tGQP4HcKhBz/2lTmRA9unbiwd5ntkh5UqhB8SK7ntYpBjUDt5DOK9kK0CgeJsqmquNFX
LqLto0opbo715o0xeWJgqqCcIPyDmx6AGuKmiDUGKUCwJkdIOy+kkb8jnCiFtRinjQp6Peq1+h80
Eh+1GkpYFVGiLR0ldMbgHjNFmB9IT+XU5WK7KmlAGgSY50dlqzUemjN1YbxEmZFDicu+trVI0LFD
SO2+2uP6u+5iXX5KJENJFFNt8eS/xGxkgIZVfn4b4APQ+JVq8RD9DGVdNloDQC+1Ku/HdMeKxsNR
WecKeh3LgmkIM2/PGznLhaRPmh17FicwXt/jdQlhlJ3sZwopmL2rFsx9cwzQlmKDS3hssYiZudfG
6gTpO6Ptb2aOOmoOlYLAVtlvD7whAZyOfF4ysk/vo/LPnw4jlTbCHeU3ovr0naUydgt/cQfjsYYP
JD6Ku5KzRjZGGyHthsnpaT9spYjMXfLvIGKY/pD4VZ3Rh7ETXEhxwdeLkFPmLmBZvSHi3R80xHeu
oeEH2tPSu9JupKfmGEM42il22c0LS8axw//C1VPqjdINIqHFoRYg3KpXyFSQcsuCuLoG7QRNnQ4v
VyvsT6IOxzc147vcaGRo3QoBws7wtnbu8gwuDgekjtfcarrIAAYZI5xPA/zIM+dv62Pq60KAwwrB
k+HiCBb5PNh+J2pvI6JSpcEZ71FaY8wuDX4aWG7u81uOg8C+3ptOBRCpcDGrWPjxMLNNBJ9CzzzB
mGJeBtPiH+effEUD24gZ+z2ljhRaswts7GqRTJg5h2XqXtQJ7HYgNfgYfj/DoraB/xrNet26wVNu
4GA6IBQij8hzPbmEaZ9YJVtrk2QL8vu5lwCATAm3Ks34DTimS8nYvOBbKkw8tSQJD8bZ4LWsTfO/
sdcUyFBqF/hxwmhoqkE785kt3ijxnbfdPGNelQ9GS3KOL9A/8B4NUmOD5NtcdM2jiSU1zL6H7L48
ITaNTv43qC0WsFIcDdL29pIjdyGNkV0kmW3jmvNqoSKQgOU/Th8I0xFZxIlv3jGQyvoQM3yDk7nE
JukeTyOu6pqquLwKNvDjm+kXKNT0AuHSz/tNcMDZduk4nh5MIffuNrvEZVnUatR8XWCampcV0iYx
6VCYPX/rTYlqBDsKWYtxy4Mn8+v2VEBbBOcWvcOdDuFrbterdyQZ970+YQTzmoyaS4i/xBro0yQB
Z1oCk7hiP/hb8Kjul9b3pSin+Z1KjglCkEN7t2AYGeuEQwoxck0t0Ei3gMBNvXtZa8Laeq0vxoi6
f7ZinqGWgtyrGEAImsR93WoFj8UoTE+9zm5HuVhZQHPF1inV6pSDqqZEIn2uH9n8A2Pv/mpzhBiB
uO9ztmePX+wiRRvvE/WaWhW938JnSanO+Z3XU1tHi9pBB2qs1pA6Z4RHd4wfFF1M6KgEOZME1EQx
UKoiuD52acgCuC6j+7mQFxhw43NoMi2pQIkY3N9103cNRDjCK1Ip2BKrBH6NaRwPUX1PJMglyEt7
BRm4K5HVPdWqHkcICxNF5u0ZjIehlS9hPRz/EzcfkKGGeJQb0FrfMucaVfLPMspK6I8awb3Z2uGl
L0hjmj66skRgC/TPZkkUhFTVTe+PduXd2D5PJ4hqdKtzm5Cw0abAE9etOhN0awro7hMteN1X+Dvj
rbf7O+Hf08ktvBQuJrpsWmYdslpr8mKjAkyNfvUZk2hZKhfGQSCOjPQj5j5XeRKG2/6yqFy63alv
6vtHcd0bPXbnNE8aVMJVoY+CikSJNNLE83Md16OcyJ7xxbzW3Rd4T9TBWRkl0zUVpW7r2by1Kc2B
k7MorMXRXfaiAoQL8l0a65F+r1EMQOIGqG/G+CBlfLBZPQg2hMgZcshW/dDN+VvIXT1Kl5bwxpYJ
9HIaqyPCKI5CWJel+Cd22WUvxUdtdihkA1wU2O6nlB9yQSGQcqqTOfawlGCaO5prGZvZ/huLYd+C
Fo6hxsiL0TRbX4j8MafdPCwXbsk7+qEkR7diJO5Grn7mO4WXCUlC12T0t1t4TcdZBubsuUSQ4Mc6
tEwDHB5Va2/BNvpHE6wGBs2oI9uOi5jWgzV2n7/QhTYMXKZIqbo95i21TxBe41wfe7wE+aSnxqIb
OaTsXeb3FI9yTl22q8vWwHQNkGoBJ/W+ukLV+qj6khUT/ulHgGchGRM2y/1yhDMDbnSRDakTR3wh
NsIL+GwZIR1E+hHBEYY4FPcEoJqxOY9p0n0QEWIPU3AySfegRmx3vWycRg3Ym5mHqaLOUlR7jm6V
HTed7DAIxJ8u3nHLKxGHzjYKxcwqskmGPLCHWg9S9Y4JbFAnPoe/yqC6eWhyOlm21fsvVz3fhfnX
1IpMxNjBm6fd/groaZoaiInACtQNhmrNZmxqyS/nMC+KaFF4HhH17ZYukmToKICmTXJCpv937SHp
2Vh0Zsvd+J1a8EXeXclWZE8ju0U95M0GePzME2JE0nRcyi3A/b0XfXo7ceAEyNE2z/m4DY0j89Np
RQTGnIAL3/3Xx/8mHBMKGj3H0bvAASel8nDt+xvFw1nsmXLK4Sw0QwkN0j8xHWt30qnRCslqEH9m
VySgromxjd0Dz0hBuT/EtPWM2hVbvmjw3p59skZZMClz/N4zX6Sv2v46KBW4eYkCNKHnkUEPj10D
IF+AJbH5hcHy8FrG3BtuLVDjEOp+VJzy4vQ43Vldbl4VcGo/949xmyeanMU3hybeV+lsUPByxOk0
3RQ0mJ4Aos2H06enVe6EdGmcGmOKcJzufnCYIThzYKr2nrN3cUmzSIvoYiMBtq8DPMd1+J8BEUvR
vVkhCE+rCTQlj+wnIDqjnWSBb2IsXH2Y2Vdpqokfx5t/ZWB1ZoAYv4MoRyqRMNRgJtr1v80+rsAp
N8FZ/to/5gPW3eGDVS8Q+ybXHrAu4Bp9K+ukOth4fHqiF2XbTAqsPFZ++be3JFTYq0HyMeXRVz0C
jCE+fcfeS9R1kEkhIFFulcFS9Pz8SpPABecKmHrx6n9irJPFsZK6+ofTijQyJ8/g/IjUX5a7ymNv
Yk9l0EbWljvw93VQ2jdTO+MgdOLYXJ7rNzg/KQ4m1Ava0O95z/HOXh3pfXKyigE3hdVU3rTRyJ12
W933qkm0FhZ3oGjm6ZHtYlH8r9rYoSCBrT/1csrEE4xrdIMG4EDy8qQhspG58pYTYqnK8LKSnqrD
byEf5vWLPUGo+knfuOHiBJ+xP4AC8XnbWRMJ7aOZ9X53wOE2IlT0YF5H+vZB/ldP9r21Yq33yPCp
CP0ptgesKi9c6O5N7O5dpXboQKb8ceZ5COiJ0cSA15TKO8VCuzL8b7+uaP9Exs6ikpy2iuK20Z99
7JaDqEtuV6mRP9u6sFCHhXCjEt/5/ZafnFXm4ChcqPPt2+Pxrc9BANlH6Tphcu+DdTVHDV5L9UF5
3aur1M5fk/S14pYPCcv+urtKbASUO8B+bKK+WGyG8aMHkZYbHum5g5c7ktnSxFEpTyqLyA7k44cx
nzQi7uDc0prpBbhVz24KpIyjRIqjv43eqOmDZg77Hkqb6lWxgcxBR99BbQAebaC59RRZxsE1fpjn
qkIKExtj6kqmAAs8mHKoAuVhZoR5Ffkl81XRNsFJNddv2osSh/iyiJf+CRBtekOsp3GYMhyDF0E8
0j6hS+7TaKtIn167DhMLGmyaTO4hgu5kxu3XDSnBYkkC4nsXmDCpyE6Y9inheoWCjXjccDibU7Dp
2oF2/fCsZYtTPCCwiGpLRdFqJuxJ4Yok+KN62lXCtkX0u6fLPlySRUvXXYCccFGlkxhg7YJv9nHa
VrY4ZH71FzUwPRxdpMTOkKWR/3+o8lwMY1o3nV0NDQqXqM1JSDJybDT6dFkz9kdw880WiH1H7rFX
loEMrVKunAFSDl1RTzEmtyx0BJsMwncQntGOiBEYy8eWB0ze+iFb4mwQ4FVFjWDqj/ohqA0Zt/wI
6YkRud/jyvvHCVJYERlhyM+0NbntSRAGHNVaOaHJiHNWYltQeV+00kkQM6ahfwy6yh7XZGjczo11
XSpIUMNTFbyVFvkhtxw/3dXWOr1hKX7TTOOVNqFopQ1JvkyQaby0pFoI747zHfu9CPuXQZ0yya0i
IDdOvGG8w9knrfY8mwWjy4rpS1LqusbR8haM05C8UNb8TvTSJee8+d48Hrn82qmRF4+RKEfn3YfX
QiUqrki9ECBY0Ohhdn4Qyt90q0pGf5hk2HyzTMu7Tac9uOjKkTVYlFW9mySRNPZtzwQgxip9T99k
bveKTbwDMRBx/L1cuhcQX2jPJAZJeunXLlogxGPzLcBu67fKNllX6SXwFZRXrYffhXQTzi46mJqj
ZJDk98eeKgqJwDrw8bWljt1KUjk6ELJzKQpdOw1xz3yyuCCrAPEAoTKkJjd03yXB+R5ziQ4lrY5v
W7ryJlcMEx2dQntb6LICc9Y5yhULiYJwx2S8zMCLZI6WEVOlHxjcEzHxdJs+ieqA5tSaXi7RkzTS
dG8VjBZ+5a+WrS80pP76ogIUS+GhhTgHR8z6wYa+xxf6VdPkHrY3phnxmM/GeClzvC1ZVwq6aruJ
4EJmdaLQw3YJjGZIPqDD1Vjrs4IvdhiA0vZm0mRWWukj6pz9U5fwJ6LUl+zxUL6u69n/s9AD2ash
g+L5aluxEOKi9CPwnESP+yrPWSI7s+L4Yex2+l9LaCM7t/NipUXq2RAhOdMxrQ8/hE5TAgJoZHmu
w3LoBkYA68VzBFu2k218bdP2UGyZz9dInSl1D8A1kO256a9RAwkbp5xnI2XL53VGtV5ykGeo653i
xCu/7eUTvCn0NFvR6CQC4d6CNGo1e51W/o6MjaG5e+YLkozI3jRvFO773OCO0RGc9NL3uZ0xtW+P
f9YgL7gLzLt5mPf2BpPmsX1rAqMoaSN9yPzdhN5kowTYPOEr9nZUV/8r3ndqVVySEdsZ7KjJNBnn
zwPHCdR/wEcLCUvT9ki+wK0OL2fQzP7pMOkNaI7ib3zhVUCik0vJ7mo3ng5mM7IIcOLwainsWylM
qtZe8bJUxY2B9Fxkc6ZNPKCk0wANKZmUaa4/54wZpyM+pxhHp5opFbtuQonG6D700tp6abmVavIz
+l2rnEhbJxbHYGp+RgXm1z9uEYKTbIE5FJBexoXrOPvSMeg7hKDI0mWvjNxZPkBkAFZiBUdLgZ2Z
1xkQN6Wvk4rfEEbN54KhcMgdJDI4mop2ZZlzN0FrueRWcyuSQBTfnvRTwcqz6nQO6vMnKOXRMSdS
PHdlZRBHEoiAx3pHmYeCdBvxws8HopKzNpANxqs9k3wwvnYPgXEKDUEapcCeGfF7jSrQdCOKGgcu
U/TVojOfDAM2ALrCEJFSR6GX8VhK4KqTafWaxTS+W9w05Bg0LQ02QwwgSuBvdQrnFfkn1zt3oQ7r
+ahNLjh/GJE2aXfOxlqaFLsH5vdiWLmB7GOHOBxm4F7+VovgB/wyE9t1gMpiaps0GRv2GvrMloJO
kfKVerHfpAE7ZfCUabFuOm9GmWp9vg8UeqaJzvzuCvhc4/bCEetZbv30LAdWyNee3UJz/0lsqpIb
JvvYlG3I5n9ik4RU0fF+Hij1LzLRvfqIKrdtIYedCd4kL8nigXlvPuQk24jtEdh1nmsg1Xgdt72H
ZbmNJA1XJe1hUCMoLXS1SbKeY+HWHvYjXRicgacvHa9ZVtRmL6nHyAQwPpGodKAI2RQgrmwxL1G4
V9popvr6Ti1un1MT3L6G9AricGm5j/Yp96TMa6uCv1WrLnyggq9PuFQcYMS+G3J8t9n/VR1fHvj4
EumRnVKpJZgSTNmqmuB+zj4jqLx3vKTAUhgU8FLDtBicGUqjjdt+hSxsskMui4ZyywKKnCS3xt0b
o+9DARzPThQgEw9s7ok8iBWUWVxEls/diyhjpM4LApWO/s0DGV4/VBKWKot8mtoj/6YXn8f+Kz1z
SVsRUVwYufswekY7w3OldsQchWySuZX9jIf+syahF2llC+BGaBhTsbh+MBZAtr8FXetDLKUXwkSw
CdYwxHAAQJXE/val67BxWeYoNgipaeTWJqBx+5N5FGqPfGY4ndFuMRcFduY7XuXIFzV/6OVHzv1j
8ZhZ3ILfL9CFWa+1o5IUNE1A15SWgHfxgmg2rKYMz80vRcBE7wfSYHHehFtcdc185WHRvtEXVoJt
Q5rXD68cLe8YtFmsQEm91vZINlET3JTOx9Oq0DFGHSp0/N8yYVubFMpWROEjlITYQinO/O4qroIb
DS8SquQ/98EezcPi+DwsN6UDPa4GSS6ja1JFJ5sHncVQ7MU1LGUyZvRdXOdF1E6EpEh7rcDoX2JH
eeMfMCtaG3ylJtiApb52Da2aOw9mUCvCROSbeS08JnO5vYKATbd/qMP5ZBwJT/y/ygzjR26JGvQs
KgY60hL9rPjPwVYJqMkmrbwViNIBbM/fWr4FE4yK4JBO9JhJFqNXLVnChU9L5ZpEqgC7cDnXHRtc
mQ8MuWnWk1ElUerzaEp2Xr4Q31ZF/5n/dAMiuORtpmy+3FyiPdstLI/mBfjATXywaHJSTPFRC2Jc
QdYp5ChRcAXgkECzm2uP0M0rKTQZxslRAOLyT4xhazZpwRxEgHIW9KdVCWF6fYSpPgewuT0mQt4o
3uKiC0s4D5hk96sy4mo0kN4QR0NvqeICACrB1NU4qnpXCHUCVA/m3SqfzqYS727MFs3O5Mw+6z/X
MLvZyowApscG4UgirXN+s5K1k1eSRHgtzo6lrrFsG5UnR0tpwpX247tffskKychgrs4UQg22/mHu
jZtAkTTEGgvWWy1eWIDarwG66ce6f8U2eTyZhmar9LqXzwtQhtcqOMRVReRhAgRAZySZ7gGwTyKY
3NusEqiGuHAiLJ/lV4UR0hP/vvmKtych0bpXXXtxMRVHKJiSBJB92S8ds+m1PjxzGO35mZJXokha
nuyOhjNz537CRiDG1t+yVBLjXW1Kv8Md76WmfjFCUDeNassq8LwcMi4P4MrcQGmD0q/3ELHx3txV
ZfgkU9Vv+PXPcPnEp/RDM2OBdIEtE91xP1qV6PTGtB63/2dCR9QNUfrxe0MjmZJQXbDmZHDrU5eC
E8iIcgXaySaSdx9FoJ6HnLYGdB9sS67FxK8qs6AW+RYtQLyQiOgWnyKz+rKU3qGin+x3CH/0ByYY
W0KUMEKcEcO20aXfa5x6hfH+NR6101zmqh0bj/Nsuio5U4Sp3MbTUIkbgqctHHQyovq+FcxiI9g4
StJT7boqb+zsbSuzKbuB/ri6nSNh6+BF7oDhAEmI1fgGllhZzxyj+Tc/RfsOXNFwfNIKdx+weoIb
VsSuoAdCee3NYlHXZQBdrLNNtVkHphuRNpqHhZtdpSqsxfDjd1Aau6oU55oKwi7DmSSbSfYJwd2A
ey3eU7tChSd2lcqgJ2Hov4l74BSBu2h6tzOCYKTxS+RJgSg/qAomzlfHXCTVPD06q7RqrS/Zdg36
fE3rd197CW1hndy6KakokrnfejoU4DdpF9s6UxTa7sJKFPr57alaI7qSGifcynhpGyUHMUEPEdEH
Yar56SuXEWmHD0AjTegL6TjkyjRtoqBnDGKc2Zx6IfSdVlBISCfgFGYF1k3mWI05Gk4OB/uykeB0
unnlJWqLEors+mWPU5T4MFa87GR8nB7GhrKle1lsEHtXzhc3XdX8hb5c6M3/wG16aNye9bl/LWXV
Pj9kZvV77bRRNp3+y80uxGJ1+1xz70hOAw8GnXjxGhZPBm4n+V1whitExl68M3Bn4afA8vEI33V+
Hhv8XISeztGrQ89AjcP0oB4k5H/CctnTW4DUlgrjc6O5xSO922IhjTgRJGeV9xcmI7KLBQYQQn+B
KWF3IVvy5h72jRdZNwszLZA16Pemw3VSSMZt4Mka5Oub7jZRLiwDxN63MeHRbKmUXKr6UtAOV2ai
ZnoDgRnmQ0OzgnrbF3CPPFDMqk0jTE6SVbo2xoUCyh0tK8pfB/8EEt0e+fUumgWVLL58qnmQEGHD
fJXE6uWZ8BSo2ErjuyeRzKwkgCW97F5SxauKErdGc7tZ3RIMMbvBBCzmdJe7o/gjgB5CotfcG3sA
1nnOLhUD90dKr2hAgNxMQ9T5hMpaSIVPMjqZldsDItO1C1ENcCsVV3vIPWnu2QY1znh5WGBPqZy9
yvWgJMslWlbTP4D5WKNjvIVOK+98DJqlEtfyFF3awsxafKENknjmdqUwT1NPXxsG9rpcjac6Lu0k
DbDEZZZ/rVq9PIxb/qjuVF8Ah5br+Vk2fao0VPmYELhKW+FbOFGXtwnuKr38gR/X7er12BoBhGJj
2DP4n7qjd1aNQb/SzmcNYBc+OGfO7Ijgxi9gKcJQWTOUiSOPSXrAGJXuevCTyN+L3C7gMV/6eaJG
strKFyZ+4iD+dZF/kaLFyuY18LiW3CUm7xpLU7PdsBVdxz1WoxPen9AW32uFdPcQJzBiiSC78BLc
ggMkpX4eYghy/hpK0/XRIQ3BP1A1S0KEgE0zGt8jntZ1GdLVzOsuuz8fDBmZ9mSloXWIenr6hGnV
NLIyWnd1Zs+fkyHx2iV6BbLfL2B+Dd0e0GZflAnDrOTHmGGwouKIPRkRGWLo+f6r3Q5PhBtwusdL
dDC8WuHDGwxJPV31tsjgAMvL04Mn1Mh3pU3VHLhZFW2SthX1ucPr/CiGYX9c4yJgmML7QEH6WO7U
4pfrnXYhD0C3oXNLsOZoCdBVkOGwPRu1/MTavk/OblIvabgYuw1rEwL35fAigBvtCAsLdqxz14bC
nwph+j0rEwUICV53ffEvG2khY9dARs1nLXPmd1D7OOGn1V9DJPnrWWGmr3mE3abbeW8FVCmaV2jd
VTqvQ/NsqSNzc9QRCQ2HKreGRfY6YyE7TZnO2/5CR75dKx8UWH8oe0Iuh582btLeBv+U4cS2RgjZ
wLmJNX/D0lkbUugFhzRjp6XfjhH7QB/Aq9WQr0GKk7OyzrKCpqv8r2nR8g+bP77YUDvoF6VWp1Je
NmMDABTfDQoA1ShXi86EOxWhK+HqznhS5ZuTLJhzt9aF2Y737imnSRfmK8AKMBJc1zw5hf5ssVyY
t6R08v+avo5tQobRQ8ZYlwCyE9bvukK8eHB8gZvJIxJhXYuX5ZthW8+yTdV5iLHC0BsklCKzAW+U
tBsVh2HAow+3z6KRDJgcGOCW4FaI/aX5wcnpxN5XsjzblkKTV8Uc4V26c9+J31wdJ4Ckq+xYo/aK
DLdC5B0rfsnEL+VT0j9bBz8PeSOBdE2zM6PXfF/aEPX8cLy8vjzg9+P2rs3IAxnX/w+UAk7JuFYu
ZLaPQlAoUbwVj1nDOqYkPOiczBYfvhjIhs1RfMyuP779KyyR6rajKgeJkGoNGRFyolXMdqwXgJLm
EuvXnQIPwR2VT6o9eHsum+W3XqF2PIxVqbFNk/NTmXuxpedsmtAKoHGe1QdW+G1Qk2Epj7XQydQl
BdCMcZX3kFfZz34cVVGnUU7Bv/JavB2n2bgA4fdPqYYxCRhr/IQaB8H1WYnT9tZGaSsYYCXLhvDt
e67W5VRHKyABuWhCk2zo6PLpARcKfvY35EjaajGUtv3TcodZOJONrKjzJsYKOgqAlxvzmVSTY7Bz
IMYTGPKC7swkPY8Mh7zXO30TXhpdpkmKHL4k1UNXnignEflJpGbAf6IOVk2r7X7+BkMPiA/5XEhY
3FBDA6xkzkdtt0Ua7WZR+OH3X7LXZecO8p1NXkq8h1C2Md3zO4TtijDFJSjcJsgrxbYi0sov6sEM
8Nk3v7zb8GnNhKpV5ZJEgi9+Zp7ITa76M56T6rrpdzN7DiouEk3PLD09Uq5xLKwYMJxWPh2W1o+8
BMLzhPBXXeLbFXv0gtLdam2JflIHNoXdwTTO1l2byf5712OM2JoGVEpNn8ECbeNZCtLQoIrlBDvD
6reeg5oVlGQ9Uk174AGUjMTOJZAEUCJJvWPp5XJvFjzQLqT9RluQZla5iSQVAdzWjLgivF1eyEjV
nUSLBJlgYxIPbfglCbJ0OoPwXCauSRXCw7gcrowa7tEMFf+P5JhuzjIiIK4woHteR5VQbK+fffln
wAFM9PppWZnsOi3wiJinVEOjrpXiBqvAzJKAn85ykZMXfERhmomiiJ06Dlc0cLo5gJ4Vqjt1rE+l
R+pRAjylCF4fn9qW50wJmAps4korU8qpkR9ktPMPd7SGibitcWLjQFSmBfR1h43GI9oKDynPKQqg
hzi+dlq3UjWKBHHZqpLv0gOOal7XAk7f3gUuEhJikbl99mZmzzEFO+ngluFSbakdB+SrWVvAWc97
C8Qu9YPaIqTo/VkRkubUaK8zMjvg+XcRtQRgNRAxKJa3I2oSGqXzbasNnXlLxFTeIhAE/Ao5IAJ4
OpckfWbnk+3UAQVmv1jomYQ+52iKr8Q+lGeekeID+nVdQdIPnMxbuvnDf8Fn7TwqL1ayRhG5Ua0w
UF031uzh9Z476NQECaNT9WitgQ7rxooj31skZS3VlAuVyRiQKzb555INXK1jw9aqixPX8LkwhVDm
Xaa4Z6v+DxiXU1FWrCPjqRoMA3E1qGbCeBncRjWKFBWBXSjjxkJ0SGOQHFBItIZjhu2NIDGIIPe6
0zIoRKwmTOxZpak+i3X86cbD/CElqPr+80Hx20TcaRUzbMhIYePwgeEUyslEwHXDra5uxQEXPIPL
xuin8HOEXppd/ceY8ah6rZn1fDu/lScZ8SnrS1Ywsta/R93reu9UrtLrFLzPGqlEzUpxymM/Sl3z
6UtHa+XsvH3YDdDz2smPIsrYSJL0Viwde0pyBdLsBC3ffOhR3Gu5zHGroDI6QDOQpMvE4Fh9vDKF
mGmA8DnSyi5bLIKapuzrm9hOAQxv+FJz/OHuaIdrS4kqcoVrhK2EGiJy17xI1aQnjNWGmQX3RZ+w
nxOWACX+TvA4jnk0vrGWYqFCHFl2G0GBuVvLSc4JwCnX1qzmGju15oD+xV6fQ265xkTw64HwlJLj
OCzu3d+k5CmpU+bz+6u88TeQqofsiBsDP+f1vPsn2Z/OCto4fqpKmu6uH2Bi8mFmhVWpShHw8PAP
FEzBfANBUZVZmnL+LcJP0yH2B6PEec9cZzlqdRu81TSXT7Cxgc1t2Qxxzydjl53c8CmWvWADjWsh
iW6cDpiQ5IZLftq7Rcl50AFDPu+FPSAqpzfj9aYxTQO4C5NTJ1IDVZbGFQGblboNxOsPGOJV5Jk3
e8CTlLVRSphtd4JOQ4oLdrI8YmdxzQYzCNbHIxniRODTSg/EEnvgo3mnXoL17aiHCjZVpiQW5EvY
MvIHOChRH2YNNiNtn4NRUENnFMWuhZyQMfVTMTY57Uwg1WIxB6Owv4SJXDDjDBds+MZMovX5xK9N
eoEWwsaszWLfh90NWYLz+/OG3mvY5akzAUGR5N/jPeoQvpZPLNzNSW4kj8/Owxqo9uJ4JLRaGREN
fYDMVaqjXiek+xrSP6UsCYpaHyjbDzph2NJn0iUBOIMskgpz6ntiAfplQtCgJ+w6GiCjNcfAoe2y
P1sv7GyEzKaJmFgtFQ0uGpEQtDViMNhVVek7gjZoljsHm2eZz2ugVMjfc4OLwe+niT0xK84nKOO4
h5ohI51YdsZUjnsGk2/0QxaBiXN9Bt/wda7IDl8sWPHe41p0oM8MfSpqAqEeuqT4VpxlbSYSKp7V
u0B/kJFS0aUX3wOFxSQvBV3972SXGHG4mjxi/Vtg0rEiwwiQnx4Tl6//ArRxaINHlIYPdnOISelJ
pvuWkd1RjIGtFZEb5LM2y7QJC59hsiKeBkcOjw+nl55+MWkKOLP0nv6E9Q+qBW+38pDDv41ITuWl
JZxaXwZMEwapJYvg+Viwp9XewZJPi9uwtOEFkajcemr6d3nSqYEdOJSjhxPUqopCvD1FDzxsHpFR
v2ig7n0iEkWZkyLDXsqgLfY3csU6WsRKjXHi6yR9hjzekhD+AQRjbMSgR/d9sBFQJiVoUZ3B/gUr
K7d2Mw5vTrbCqZRaXr472DsaQ1OmwHhdmsvvwGrM/OnaXo/Eg5Iq4RseO/RtQi9uoAs1wk116SxN
aTlr76pgoB/nqRhIXt/t9+TOS8K4uGjhF2EM8Bk68U8G6cJ2Dd8JC2Amh9SLmI0ViQouttvNX/z4
mP0ENMvoTqKJ1XYpFdAvPRStSPp6nYyAA4sKXcazW8Gd7GeJ08qm6fb7ctVN4cTEhP4U4dihTnLq
deW0y24XcpJYc+ODaYLCCrV7WArct6ft9FWpki5O/i0lYlWVJLtosp67FSCso6hsj1H+nQ3p71wm
EtNzdV1pHo5N0h7E1xccIzD8j1Z+8OgurNIUyo9/eGGD4gVJlewTZBZs3N/BCT6EXqjLq53JlO5q
WiGdGf3mWMl4KkSpS44wuahJTx+RgsInZY/kWViYuxaomzA8JbfjXCIJH2lqyBarFZ1XGX23nKBr
42SJQNGobLc50OvW2iHHqz7k1FWxck1nbbJxERYU0aTwBfb8JfGa+q7FFJZrQJE101Lux1VZ86hI
YaFudxFXIXQT9ecWwgSYYM8hDN3YrYQLbqfNNk03/4brEXkCi9JJ0Qrog4if+NSA6b5KANtb0k8T
jIfgSpmK3ztnLJDbznEOdEYSFncG6W3f3q1T7OdEO07mxd/pyuyHEoUnczPLISYcie/S4s/u+fLy
b+9fnWDpJTdI38LmDUY6dyKK8puiBUY7LZJ+JlwFs+vyXGo8dyXnyKQg+6ZbToH9wJ5X1Ck5U2mN
+jwhfRxHACJcarg2Q21/0qfVAEhMVbUuGQdZbek0kqgWvTLh0Q8xe51ulntnXifICqqtQGP1LKsp
Bdyok/yUPEPDGMeWOPJHbD38nfKU2Ytx/kf5R3awomXgnnlRDvj9X74E5khvo0yPFfRLvG0kNhWQ
0Wfh1ToJqCoi6vzCBZSeUBLEKiTmElqzUevvtJHO8ggE6vpwDhOUUCtyrGwBBNQ8owRLOsiQufjG
8Rify8qv1G5ghV629DMXLYztx9SzsEcjrvq+gE82Jhi4O7b8INrq2fyscTK7q20KzEpOl2gxgYuw
nl1lbCyB5fyI31/x4J4N8Ok7iZeF0grCTPHTx9+5C/3f1e2M6yjeDR9AunfWBvhBF/16IpXn3ri7
DYB4OwM806xfh6zhwZy4ezXdbUmoYmSwpfMHdv+QNnhwIHkJTqXmSGeDDhDVLd5OWs8yWyjD90Ck
c81otQvF0KsfX8ltmU+qEZNn2saI6r+5BV/EfVRTr3TrzD6lRZ118zILq9mZoV2nzQpZI4fX+D3b
w7rzdtizhLkqE0v7YKCn1g4qd02Sj/hGAQx5+93P1QTTWvMJ6YqXeR8uInzppwaLkuXkV36O+jDd
6E0S5HJ9x0197zWkXDyNHWU+LTCTExS7Ht7pv+T9axew79I2NU8uf+XfUnoweG95XC3yD7abKsVe
zHNIqrXWa9s5DoCVoP7W1NSrPMPlzyzmaV3qPw0kDMcZdTfC2XjZonYi61yjQD/Nq6I5OK5JICI7
lgKCSHVbp+GLLa/gnH1jMD+H3WbeuavX/v6woGR3e+nqgupgL2gQdqtPzn21y8C39uSmjj5yX5SD
6Tj5E/G77SeK0fteCQO/XXY0gSpE3q0JFExGe5niByXiCiuHGaHMhoB4Q4OmfKdlYTgHyv0IphRD
nysntMdaParlQE+prDVd2fFprHldts2kJYy6m642pk7Ojx9N6Ha3h72hW1J67Ear/b2Xkui5JFne
4zBuF6X2Jqxb8QGZjM7xymvo+jzWNGdmpBr2oMJhrW08AeOE/m9qEBklnvLqI7VNxOCX0c7U/lT2
fI+PSOdiiByD1rs/C0zcNC5L5Ok941Y/vngqkR14o6VrXmhsvL6veu1tNV3Siip7mWntaEUxlU4k
T6QOi6ru1Tm7p7krWqzn63dpyIf7WmdErbIa6czcMP2+3FNJmiM6sIfNjzduCsEl1UV1a0GO2d67
9j3pLby2thBt8Y0B/ZuvEdaLqJaZWVtfawJGFCvSSMF9ylUoPYkW/fmv1T06/U6TwQo5vQmJhNcG
LL77DqVk7KACHxsoTF+0VnZcSpAwYrgP3MUTmBT2CfELtl9JFVLeAfeud8z3+RB6STd9WwiVwBaY
khgEs5n4LuVdAlU1bWKCw+Z9hGbEjxIcrA/UA6rMZAvZBVtaruB7LGEFzKgcjNoJbM24CasexxMH
dkBAv3dt1bhAttNqaWKmmVk0Up72F3LWCsWBjE40faNJJvl1tFZx620gqMTlKqcegjNWqDpSixdE
KdpKh3fS1R+dsIxLzrpus+sNMgjLwUcI9Oe2Y2olbTExUaAwP1w1qhuETFJN0Un93AnrWvSJjHHx
4P5pembo+foYGOoDV/E/HR3aKKgesgVBiZ6tl9oA5lkmTkyUc92TNABeHBEfUWvx3BC02NuNqmSe
CDz5PU9cN38GROTLRXhHxmTo8DXil3DzLV0cWLqthJo3AGAXyl9g2asBRObkmeRZEX4cl0a30Isy
sLTY8jtqh3+HYyPV4xAFkYP8sZ5/QrIaVDbuKRpICm/zdSXCCGnWpbZ5DotQ8Wz8xWO9farBdB8P
ASvV4nbwpGvcUFgX6YhMA0H0FSxJMSPqoFl1G/4H7tSpQTXpCPEHzVYc+Hq/EmU0Uln9jxmIgmxR
uJeZK1SLjI2zjCoMldduXif9OSY4XB8RkRI1im5ZwZkF2XEqIyHZr3ylERzx2F164GsHJloxOmNn
uL3HoY6Z5cNYmW4M9zYykjfg6ZsVFaIa2w5wHfzvEB9vBu4eXMUbgVTEws137wjYeZY6r6RVjzL4
RjEBTc6mYFuWiug1yQDF8ULlMCp2eq6sNAAJDSorWOC3DPlH91pYoqNkyKtw5c8WjNsmLhWQ6Ydn
nJScdWwfHpWeWFm9d1mCshTUykss6czUZHn+cpGrFwhFup4vqABBN5yr6bsuJTIehy2dBdF9GBhn
zMQY8/50R1cu6eCkVH3I5eDnmR4twUVK++I84/+6CYh9wD8/K/M057ixpQg6Cdxp5VwkPJ/kqvid
VQ6dngnByoiEVbXlAGVquxEi9JIcyVAknpom7byUeb4sH9Xwm1Bj/Ytene/43fuqTF3NA9164cKP
wZbENLI2mXbcLHJaGvKclBA9YAhM1slF7T/fCpaybQpZ7848AxIKTcZHcm3IyQ9hJYb9zHEQqYhn
a7rAX3Es2G3QfB/esMzjZCVPTIniq0eSDYaga8hnG1/pqUcry7n4bokpdLbpFQocooIsR/bYS8en
4kV+K02RD833CvHpNGe3dXOKTBEoh3YgYICNUxNmO4louAidWmd5LjkzQJFDuakX0iLIrJ+aeQYe
BL6HjDnnHCYJrdlbStr2LhPDJMWliffsslooF2Nw23xhgWySbc3KKHq3W8aDEPdaSD92EGiGbDjO
5LplWl4aHfPagOO2HEN+t/VRIpTROLNOWeVDoOCqi2Btyb5TnnK+i2wH8GcpA9MsoxEG4EPoKy57
BK8a1vZLsGkWx+piBb3sRJjjAiGMdwkQL2CUcdKDwSKpkpm1k7kdRyfThRBwtiQ3j+iFy77H8/nL
WqJK+M7CYc1o/sgyC4mZXPbLwYPS4xO3+9Hq4n2rV9rfEpOcJ78xJjZws3rPnBg9pBWUqyXwwIzk
o8YKLWmJ9dNcew5HqzOYlcnrEhPnhJ+MK+oLDfEr50TM2hw1IWWAKYr0gEMHyuYe7zSFaAB09N3L
jSEuahIcwlzKWtdE8KcowfrLhiSIcPj/4r2XdsXD3Y+2FwNX62krZ2hvIDD52d5XwtRZbkowWxMJ
bUgilerHqS5YnmsaAxyoIxE+fGKr9QWrdVHYdV/KtBZIprwW1EEAdHZ/3iMJoVcEu587I3mVg3eX
0SaROGgioCAKvVs3VpzVBNPl00ZRVAogXV9jexZU+3NAj/MOhj7pIdKyQjT9JbblwBgjCjJX12hT
TSZ40YUSTqI+pjCEhccELxyWGQIJWqGbNmJ/mn6xaISUYC0eDTSGxAq1EGOqWhJIhG/Z7KsRudfX
7JEf7LySB19GMVkxkgX1eCJEPr9JoGQSPDrqAg9P0aBoK2pC/b5vPea4VLL3knTP+9IaoPhyJKyo
6uIOwIbamxxNTvlFTuXc5DoZVoNi8RrqvD6HUPqgSOp6mXfsiikC95WyRELnqeYNqBe24I3DPqZ1
+I4L5HkdB80ccdwH5KxrddigsiPAbroWUpDEAQ435805VI+BGqdF7hc35ShUHQ2luO6RII2wolxQ
V/o0D/ffbylQiUk+mbqH6MFHGvtBFNM2uIO0uYNJ+/6mNys+Z8CoAQXtypI1fABIuvWAkQDdAK6U
BIWbsHue1lPselv70fQpmAwCDVgVUH8LCUlKH6JVr8hHmpDGHsh7QV3P+0leAvAFI0/ulVOosJ8c
mMLCUZahrPaZOWnwi3lUM3AV5JVJ28LOe7N2qwfvMfmRipvlcL+0MQhMvcOrwAkjJXIkus6wgMkX
yaWxUvoRsTOUyQN0EDtJ/fhgIFk2l0uborV0fj/bzz7+urt7ZFl+tPEenK8DygqAou4MASlPBGKS
YNnoc1qhNxBRr1NS6fszMdU8pNaG+Y36YsWDdtb4WHsqIgqOH2HefcieADyWE8Ukq3+b6QjTWADp
lWAMVGByuKYxSd8xEuyI3FiUy0Egw/aOgTqDFxVx5kJfP21Ry7ZsIN0+/2+M4Vw9yR/dW2zAJZ49
lR34DzxY5jPeBqFNIgL7Jjfn4BnmTsGjDn0iwxnqVoD8iGee+rGic0zg+gFCSzSs9ZzlLYvJGZBC
WWVXqPwXg9SK4wuenT5A0o4lbZwx7mwAErvfIqjbQET3r5baMQMY/bWoVZ6Ed5mlgWESPR5PQLFx
IZAqLS/44VcXjN9j8l+rusShYidbup82qXqp2pRKectpp013+c6G65hS9khRNvBCw1dbHd0Sv2oU
lAlaNHSIUsj5WS+RAnRBeuN8ndZNh3/fMREbaLQrutKD7e3ae8tDizUxCel77plL/DJkP+G2ZB6L
nXsb5XvdJa0ogP1BzOIwbaDzlDlIBPE3O5jMNR7w/UlrSjlAnDTm/YgbqoRWhGedj1VvxSyumcsT
E147MEi5JfOAUcL9sIZF4LzEvA8D3O3Y/wVzR1KKRXQNMGkPBTBgOUdNmmkEmdMJmeIgyF+tlwww
OoYOsVxuHT+nT5uKhCGiQ/Ire4FbZlOkfhZo6hWlWjf6N0d9sxn5m/ri6vDJq5573N9++OjVjH7e
iOPozY4Tf/bRxUqJJhYKNLhzJasmXnNVnfRLlhhQj+55oqZeGB3pwuFVl/RK4FJyL1XzVD3axUpA
9zOzz6kLEV28Bv6YDrwmOV9G8v4FSS9oVG3U16r8HJn81IOqw8WyS57uf7x3iILdLNDdTFuLYOFn
gpT8vNRbW+MP6peboWj+V5KYklCSveHAGOjvVv1lZqidn21fg2xAuGUsJBdzBcu2JAY6tNw0Yqls
2wHNk9bUuXrG+sbsaRdqRnzxX0tumLPTnDQCCfT3tSXQK99YZ4QsknN3lz7Vl5z1ih3rQXgV8zBs
rerHFIfVbPKw9xRWXAQtU0H6ZUiIMIXbA97+dJ+9mIWzv2ZAPfCj13paQi24AxCObCHlBp7Wh1HU
ZZlrLJvwYsLqMeeJCGNQVHms+3tjUxSUfEsQTyqewJBO68e54Zh/ROwGmORPfa4zOPfsCnRwZ5zE
tTs3phL65FQh+39fY2x+rDDKPJeSbKrLXBC1BOkgQJHqzhNe98d89O07f+lx5oAEdidO5DEy2EUV
141Ej3cVhLGgxUFvqSeEx0laq/VUQ/P66kv39S/O92kNGMmNR3F8/21BvXbHzNcbKjV+ETVaWYCG
4LIcVl9Acbhjia2XREWa4wnXKcAgMqprcLKeVKqn+v86S2r8VViy+nnQevF8+saERjG+sf8wlDCb
xpszQA4Qki+spXZKPZiubTCEEN8U1PEk3mjVJ22i7ziVsjJU0/L/LX3jo7tCXudL9eDsDNCuDT+U
iJ4seOdhdwniRRfKn+wPnHWd+qtyFAzxcXQ55NFn63eFWmnqjm6cS9gmkbTyeXRoUlKS8j8kW4RO
y6tA9kR/Zu3cgmD2kgV/Cb6VC8GBKca2kyt0lCajeRI2QMugynzx3Natl69BNwWVDmxm312neCvg
BOa2LlwL/RBga61aYp4bXvIFo8NgiR1t/aF6W6KU8HGl1XQ3WgIvwj5HAXUARLZFTI+W428EDqdN
EJgrs9ztCQejJ2z0xxSY0ZS3m892uyZBRgbDOuiIqQOSjSWtGodXSCZzowpWM6PB3Ypes6aoXfr2
DRq4oojIv/us+nszenFhVYBKWMaRCrw4zxtFc10YgRMEDHk8vCJFE230FDUbBI38BtckEbSxmxl7
NZbWpMsf1zOdRQEEtdTYYGjVvTDOsRyvWwYSshGT8Q0F+O3YAAtGpoDrQEZ9BiNwo/SoTc0kZccV
o00oaruAnHF3XuizzxVdcmh+krnNmG8apYErvJ/ptAFeqWxKe+hXfo41SWQnZw2n6LMzUrvQSLgO
CurPhP2SJhaITM90eNgjCTlflUW0Kt1DkMamc9/u3w2BBQuwqYpp2vDukpRLqIPsBWrEuAglSHBU
dZFkBsvgVHLZEZN30wPQxQ2BgTb5Cq5dbUXoNgkSq0orP83jYXMmvQOZ73h6NKRfwg7fxzaVGDj7
glQzcnHKZp5ETlP5lTGC5M3PVSgKzDpx0/nSeYelJMNi1OcocmIY8T9i6yUlgSVz29/054IijHzb
3+lFYNQNhzp+z8Rfe0bIHLjECR1KGFN5hwt8ui6h14BVXp8t4zDNOF4aHArODbiUNQ51wvmTA4nt
kGXcW4hsuEWnDLlQWMmONkH+HYi1AinRdzJl5LIbGmEW/NrATe5t5BleTDNOj4tKG5fchsiM8dtS
8zHsh4s/MueEOUr7w5E7SgGV7ixay6ncXkGWBGqnoVnlq737rgkpXOQEIh8Vhk4E7DSbijD5U0Bo
Q/mAq/k62C3Eb/sCM1e1tzD+VW/Aa8e5pEbQbWZsXHv/9ts2B37Wx9xmqodb+jqT063nRIK1yrLa
cN1aH6jNYM+t8AaeTqNoOmvesTzuirUgWJTi4Drxk1jwthgQOajNNF80HOloQGYaY1n66HWa124n
Dhp7V2WPePFOUlO16n1sr+CM4RSnwZzRPuS3diObF5MNiukexowzWsqnGiBu1V1HX/SVK3U4/nye
ZF5Gy05AgfnrtCMh44pqrjqb7jdpzu3Gh0UF+Ix1UMtSEhZYYtrnRHEI67LA1Pj2BKosikSJOtLn
zCOxRIqTjgsY20VqzBwPSDFpeNjQuk81dudPUukK+ImU8o7YQgB/08k7iGUa3WfOXeJLFF9K58Dm
xO0Crrt3mdElWcWssP0BwROU7N35kHc1Wsbkp0+eAckXU4/2Va2PKBLPYzVUlsX4cdZnX10MAB2o
vok5CTgLenUWfZg59MgjVnlCpG6VvKFBqD0vriMtiV7WeNoI/+uYJ/d8U6ZdR3NvmshcewYbmCog
TSKONIXZ4Fqmyb6RSd8a+udjb832WqX/N6KYKceuWU47PYCrXHt3XXecw5gM93AfdD26DNTDFXEd
V5mraSOd+3pWPn9+9z9H5DSqyLt48uPCIEQpDpyySfuTcIxfTCcYf95Hv6L4BY+tODIHa1kTwmXt
5Fcv/qECDsNXKH8CxC6pteA/xcsdeI6Q24kTG6Iq+u7JpU5glMP/Lcp/PpDftOxRMs/uCzhft5om
I2p3/ixe46Z0t3DOHsQM4wnDW2/GwBQrs5HE6ZcxemozrLAh8DG9A6dAdfbuvsrPCnTDg5mnW97s
OmY/+9GcKtNho0+lhbatEYHNwEhK/8ibvpASm1rGPH1ddWxcJb1VJ1BYVfC6II7hWaid3kaP/IMp
3ITfefTescMpXBE6NBvqESA/RntUYNPuGa7+5pVXgzBShZLm8fusC/qpkAwQFiXAPsx/z9wn30aX
rBddDTuGdX/a608wBZah7/ZamKTuGDPLozcuydFO/sYQd7WsuVMFdwCBWQMWOV+R37XDOOJehEAG
f4VHq5xEk5focYrYPhCAA5NizOOlGQTk/NAMwSnzftjCftEAEaEG2hZb31BTA9o8W/SiBQD+vREP
yT0zWuuDx8+bW2LzNIaPYOVV1QokDkmtGumnKGsXqtYI8GMXXAbzGVlgPBgLg/dNwIMbWl6N6xxU
ug0LccnsqK2cbHh38+xDDF0O0JyaHnerJVIldp82/i5N9LvKWQSTIB02/xMaOkMtauIWmfIKyC2B
UCEdVn8YLUxSmReo1EUmhjcjMZ7cVInUcTG6nLidd6Iu0vrF/cZ+5Qw/n+RkjXVBZcS3yOBt7zPr
tQd7V+H361lwVQd97HSTzml6OLx07TIcEiG6VCeG6ZEHi1iMNxNUK0ppQG7Q+29ouV8E/IYXOHT+
1P3fQQfROSahfQVkZ7DFKlf/op3fTN2d96L+/YhiTAG6WNKHKh0Lfz70llKAkhgJlWx05hb9VOqY
Q+R0Gh1sh0b4/HWoJ2r5BppGIDALMKYZ0scFo0Y2aroXpzaHTYiF0pXWdzTSHCxbjDftXn68bWxJ
whm2rIU86OJsyCpbdA+4cL5rpVXVyxgOsZ4rMKWJsswcfGTp5sag1/WU0c95DFrLd+xjXPxujuON
blLc576hyMMFCpN1JmazefUt60/VQzgzi/C9URUBLb/mWpHR9ld/xrxCt3qmdWfnKPD30mD7cfO7
qC8oDxMOJWe5LdAPJelkL5LkxDyACPBML4iVsP+DVLRyqRj7GNVTEFZW10HByMzV+skCcR/eOamX
mB5YvM9gqxtpHaO3FQqal3NIPdcNlg/69uFfl3meAs9kzegGTqf8QxNgHnyihK71HI7ZgzDxbz5I
e9vtbzRURox7EKXi4tt858U6D2HxBFPN1eaNDz7A0Z8GFdiaEoNOz7aaW2w2qBKnnsqTDjpVvWXh
EiSG9UFoo0uKjUA68HjRH829m/eXJSLT3MTDClox24AuunOhsZASZQ9GrWO/X7LSwZHzVfchJyxn
23kg3HRdwC92SZhmHzqQrp6MUPUwntg659VccJiaAPFKWXsUumNFV/OXXsTjiB4eRVMJT+H5EieN
Iu/rrrfoEt/kSQvvfS43L3775dnq3Et8tEt6ANoaCT4uGue8FRibSoaGQqzT9wIfYCVxTT0PQLU8
3oXsNePepaaEzcQQLk7KDi+UVX2+hT16nLUrd/k6L5kpN2K6LvA1+lIAsrE2y6yP2A6s2dxfGvbt
74BCK8OtrhX6oKW2UBLyl5Abw4EPcWKie6WXK3+4DDia//kd5DTHZd4IDZoaEsGIcbHlaOd8y/iz
WsMZ+IFGJ+z+MhJ8HeBf9W31KUMU81eEhwKeyugEoiQPr8l2BqFGQyFJaO8aFA5QNDBlQ6tAF9iH
r9fQyTa4xisXizUtCba7qcZk1mMG6ZPPNPqmKJr6Zl+zlZdClR8Z6aS4LSZnWnBemoNBd+WSTjp1
n+BSDTsPRwKa/41P2rjod5MW2KYXzm4I3oG6jO1tdCBz9VCg//vKfiXAydp4WZdW7v97nioMGMTH
5lJT777oOVpWZGlLJqQu2cMNKPGUw0SBA5krhGwU1TzTzZvSPWp85IFSZ92vLZ5JWzfJOeCHBFV8
pYm3arR7f4BcsiiNvowAuRKZsXjVgLRjLdW5GtDPSGn/QGdKRE8E2FPmsAJ3IKyA3niPGNNs07mc
kXlZbFYx8gpdjuLZjKIqXChj+Fk2YEiuvbS2Fu+kCxF3tHaZ/5NqM4kYdvLZjKbbcbRvZWdQlkcK
jfUxoEdzlrr5K8BdY/4Iog5mlDlkJPdc1ZmdJo5rwjwfIt/xxY3S8/L+uizEC5hvb85QBvy8zwco
IRo5yubnlYy/Kid8PU8XGBVVaT1MhGln2BUckQgkG5rq70/QT/uwvv+0hfVnRlrIKUiKvUA578pM
ovMj69jN/wGlvOfxYFQTjsaMb/22j4ZZj/RuidOP4ha7BHPzZ8rn9pZOtjJUjapaB0aqCZtwiciW
HFHcA6cGxtCY4BJaaG/Dmi3sh6+HNLbA//xp2CtR4bedukEhUaN7yLUFyFBxBpMXeLCFgyDtPfnM
epVrbpByXT2udut55xuwXM2UDJcY8FlJzlpcvCAnNKSkA2eYTd307oQ+mfMD3DODI1EOCf7A7pLA
EFy+twuzrVfEU2zymPJbEkqRILR+OlXjXP5TeZIz7GIpawcngB6H4RDLMbvwB1RhwVlLlcijTEvy
BIjotF3/Q6Kvi9RNmTNabwM0RiGjak1SQ1AQ8s3KN7z9l2JRTMZYuo3oPQU2ga+DZvrFzMRRVVzx
onVjROrrMIPGEKu2AHzrgh60bkuahCoNj4oozi9sySrRfdWP2P82R90jzxfrR8DIhqIJPyYUSV3u
kLuE+SgAGe49p1In5T1kV0v6dxZlSrANk0547Tga/kkne06IlT1DUo9LNFU6WAm6Bp/UrTECOZ9u
GR7Vw0+s4zqXROKHddBbVVOdL3/P5ku5gms8ggeqvIbNXuG3kPgU3ummS9HZGrdnnGx9DawGGFbw
qmcz8KC0ntuz3tx+Qqt1cXdo742Y29RPAv75qgdDkrnYYDCCIzWNoOWFAkOLzxrzFnT+LhEqCcXm
DbDWNNJHZyF7x3Ne/waNIeR9FE0H78PBvXkxZqIN9NW9BtHvSTiwhjJBOyHcFNWnHxciZJxNa8KY
rwvuRanP3NkGUzsUFZW4SaSPHUJ9w412rrd1uDyxM8CpwbvQI05EXUo96up/763hIFEYTYLFn1Nr
L4Dm8a7nr9H8BpqKSJ9KGUUnuzW5BaDww52nrmzu04txh0Pl/vmUNEwRMxgJ4C3HiZJiF0jMyEub
3blh2Duk4Oz0alGQefzHtpKBVuFRC3r3jZVE6gR8xxF+Vb0Hquyx9llpYfqJpO49lr/v0YG8JKBW
tk+RGMy0MA19+HzCOf1Rg5MdgqjFqCj7OdgKVAnG0yPT/KEvUz54upqUNs6/k45C3V2uDTD+LQCF
e7xwXdOGJhsUn3QS/Kada21ksocPtGe6JTf1bRwbMf/+m8uw7T35bbIYB6xVjOTd6G3cGE4SNBUw
a1vKdF2xCaomQyZ4Grzi6S7rqLvoiXNktKgLrLrfSwLEKLXTSsF92i9WdBbKrFpGdcjFF6Io2qOj
sN4ne8hh9pi51pC6c48jGwP7OYt//u5ZDuMCdFdOd+G4Ew/ukjihd+S5kqDAP1RjrGwU3RoqHOFN
WxfN2VZtaly/lc1sXNLzGZD/8vbf6UXfFTt0J5Dj8tw01JyxPqWquMmVlXH3p+MByNyGaAgtfy4w
QQYafRF0k0hclDl8k7Th6OIOIpn28IGKMm8UCUr+sE/mY0NPDUBS4H4/89M5a1U/UvTdFP1rNWv5
UMgKy3ZHk4okrm2ntvx3WyBAo6XUP5+wlIHOQn0wXhFj+iV7PBYdPQbDXZfW2AwdcPDcGYV3doLm
YxXfojU9gq3FqAPUAHbSMJO8uubrICQMnrCkABt7xK6zRMBs9z1TkiMXouY80UOgwviA789p6Bln
cFGldKEKKIZ3PQvBhgQw+RuPS/s6/SwjmH7gvUDT0nOkOhs57aTTmCyCc7xyRZoKgP+bpYakXTSg
uBEWiGzv4OhnyMjLFRn+PMk3tpGOFQJPp8oXWbAigqznFrbDK99v9pG3rcwEDMp1E8NdXJrB+GmW
J1Ir8TEBWbeWVQCsyC1P/l2SIhbaiqSVuYOzDAv1EJGKY1cM6N8/sw3FUrQapJVomoEBK5sv648o
EEUUBLxTofNlCjxE4T2YWKH68C/gTeX2GjRPFHhT5hBOLfsyb61+BL/m4t/L2Rw1oe3qU5koltlo
Q8JObqBRbh49cqbqYQQixsK5gi7Oe7byRYjHR655iV4rhJCF8aMjMD+ggJcOeg7ZXma08o96GK0o
C84fuAFOhZLC/W0wAuq1fRjyzgPzYtPR6EZq9R/5nICBoFnr6r/YbwgJ6YKfAkLkWoLvSkWtyl8R
QOPFhBAGJS/ckOaVSiL/T5dxW8mR91QV63ERL5bMf5Cr+od/c01OwEn9Q6ZDNK60SysuhilOtQjM
lYKndyTocqT4qxdxQ5ciVNv2XcKprDT0yanDo7zqzKaUEH5xyjvag7Bcu6D5qc3Ip+Nbmv/yO//v
zWJHUEnAxLx/dMQ07cZ7uwXc7jZXv9pjX4Z9O1DZ05/hRyBih6erheis6hO/1K0Ui/52qdBPBIAl
Z4OGgVEgR2+l15rL23EZR+QqwopmZK9ev5xNA5o5Q3fRD46tjNsy4FUbkvm4ckfyXncFRukiYg23
LUtT9KCoOsBUS7XmM3gxVcy4x/N3SlX/BFf+vVs+bGkgf9dpSvw5Su/+Dp0+gPJ8O4uyTmipI5SF
6hAePPYRuyl6MaF8MJyJwUb6c1jGDh62evhnmE04WyuNMcQvkBBrFMx55olY7rGDdKh33o8CbSrm
iejgsC+K5K9yYc4CvvvkyNE9YDZ6GvdQb3kg6lU1mQy9frKk9kaSXdnkRyrqIE9eT8hrf0jSld5A
jnxg4HZ+44AO3MMvnqJUancEU3n/MfsXgfQLPEvOtIOmRlhtiffD9gfSalVKub66dyquJIau5Hmd
3MNt3VlwMDKP4vsrTCqZ786swqkC1cwdw9VUlPYw/2p27b9zwI/RK1/t6HQjNFZkuZvO29PQVQLz
kkX7eCTR1jvSzouA4nsHEOHCjaEaU5fc6RVgX/ZSqk9eHZIoKa3UslrTNdSSNGfnhN8fVrcSHiMk
Yd6a0cjt560OWJdGantY2O/FxEs1DLkNr9/L+NuFwfgwt4axpvswNQoNc3cdVnzLDp1WIFiOdCyL
mx5XZ/IkztbtJkVxj2vMiAjV5ImKmTFNOSlmvCzK5rcj3SBXVpf6RLma+a4acMAkW9noTGCr+8Dk
TxZqJcHbS75SuJkppDmWUNTdtxwT/QtLmIaP/nhgxazyiuxufOAzFjyH4Z/zbNsWvCzL/qHkHPIE
W2HoRV+yZ4dVEKsHZl4GaRy5qfLgVgWGNVgyr4Xu8NAkU5LIFBuRnSPwsf5LiLOl368jIJnDtQwg
UuNsvvU4FKXfVZWIXZ6QZm5nOoD0ff4V6GCIvqR7ePB9nrZ6qd3LQBLCmADvAZwYYjvsf/53JlTp
oQAQ9NeuSaUaqB0m68SWMA4ZzXWdHnhEBqDWMf9sqKxeedw0ot1dRgmteW161QAICaIKBU26OSgX
1geNn4oiEEZyt9vck0y73qb9tujiooZHyZRaJ18TwWGLVnBLlT1t8LNsIu2nWB6kvKuwXkQdjrlV
DSjr0mQBfrlPeQeTslKEpXAR+6KOsObrjeHL7EvYtRBOrdeKUI5d0djNYYSe7+oN4PRWXBDu2tFk
u5AFzDNSRUPI0xyyGLzKSe5v5sTm89xeq3JR73kS/boF+cxYX0yv5tunSnS+9ExmqAUxPWeFXxtx
a4WQMWHTQdDMp66bTlF0Qr9e7rCWnfMVGZ4Ieg21L7TP5qN9pIWn7EJpziMil/vXDbaUF/M2Ckqa
castxiiJTVHysCghl69H0I5tSOlNkdLdpEt8KiK7FZsEQURl0WQ3wXGQCKUJ8w7LrPtAFMju5Lik
LiQUwTTRxUT9oVEg7VlsXEkDYXYmzTwjqHdfhSgzAq2yrT2wgx7oPfyA7rUhHOeSgP5Wu5KufaSh
4GDMvbFtdQm/hnRS7LNYtAqld8gpU0b3ewqp1za04LMMRp3BCIQAOxwitSCujtmlJ8X/L0vFcLO4
xcGHt+JfzjProQVU+xY+DHU0QlHj2A8ba5KoDvCc1Uxw7sB0yMzbuVP3e22igtupzeZdgHJo5QRu
zqv73Lj90x/4+O7TRSw8nALNx5A5FDGtAgy9q3o1TYO19jSHWhilz3sHIBqMgU1TNGRazKNEaaGw
nHhjkdKjkCh9cAbNDWh0zweVvW52fIets3lyXVsf0Puakpdm56yhSNPrA6a/Ozqy8clT8XqVIyTg
DYGbDtXQ4aGwqUXnxl4wrgaWqBBxX4OXOkZnLcx5YyscVBygc81cMRG46qqunysitJ06bk7XxDsH
RWw3NRiCnoRybksNza1lSN70M6NsLOOmNIrtfttYkbESAjFxrwmro1ViDTjTC5kf3wje6uuqqOnC
Fjt7ORyUaUDEtqU2HV66dDkjGrpphSuaYqT3YJ82ahpdmNxHCNYxV675wJxEfKs4/ss8gBMHP9rA
7khBBSWmSlIoIEBbFSE8gutGz2P9ahVLhhqxg6zxmwy7jH8fckP4DJr7k5jgDN/voauq6BRwXw23
PvqJpvoWlBDBdkRE5OidwXg7YYQT2zEq8unLZP/CD/NtT94mbcbIuzyEnMKycwIG0ktl9eIIDzej
DbH6lVIjphqOD32T5ckqoRZITSTzTNFcXuhEXXkqvoRhJDXfDnq22ctZo3hxXF6I2K/gL9yzZb2p
9vG+Na/5VQanHNBPyAbvKL5ZaJUQYgGKLzuPZEWB0JcsWTyQYcc1Us1A9pXVM2DAnS4gyXWP/yt6
+td57wwH2GB2oMwd9Liabw5z5bUk0dCHAbcsbllXVGMhyNjrxfduZV9ECf9chpYWqsTtxqdAm6D5
IccNwKkYnxU0Y3ICx2jhIeqcDx9NDKrcV5UlwEfMtWTUDD7IdlbcgrZfjWmgiH8dg6W6kDpLuMYo
9yYZB5sldCMfGdTkCm3cyHT5bEvGSdg5gVtU3v03CXECzi5FHX7OJImLC3vMIxIn2o/G9Hr7mEij
oohZx+rQCLizNkNPdV6o1zfOyuEFPWLdGjM51u9qmtjtxRmo72aQpIvMjH6EusnX43XetFxfrHaM
gZdlrx8YEVkCQt+pL16kXbyjtmKX4A1BOda57bIjFyTa0cX/roYRRqnAo2KZlxXLPp/CYBTQx0i1
E/k8F/sxsUzfv177dtuJAtucbQuehGrkX7KK0IYzBoNrujx8Ic8DFItaqgG7ZUuzNjCn+v2U43j1
FYNub6BHeg4wC9xrA2wgzXZ4wNSTkhRZPGqgSsEqwVlJH80hNLnODBWlrYUgG0lbuOmn2bQbFTfc
dP3GwyhrgSaUJW/4xMwGvCKLhCGsDcPlLB4F6cEYR+YygKpGFhGKR5Jq/KtMD7sTfEj4v9dwYvpS
yse+DiOkkIPefvfSe1+4Qe31YpG5tvIGUiymia5eU/vPLB1rLPry0WFU/DofCeO72INahHgvBSrf
2c9nb600RLAOxRLLakEss1j4DmOY3OyzDiDZ3w1kGTj6zdsksTCgp1axEVwlJ4T4xdMR3LEJdmXm
WAxuoNAsA2QbMexV34ZqarSyhIIXZPOFjbE+UhkfR3ilvCzeUk/3l3FSPD5iE6mDl3eJyHcg7Kds
ISHjTSEyluFVFpi6hNB/JN2/h+X9Ds+JfSuBNT5s03vzcAcCIW67OEoVqxXpXpf5SrrnoIggVxPJ
w8esgzoL8/JVK23mJecdBBfxg7kbpfNdJ3HLddDGG0yFfY1wbpqdNyVjfnrD10icaqUCow56WNOl
ExWnxjDdnIJbJ2QtYeE7NtL6z6KKuQoKJa/iX6zsYU9yKMkTa+QMENVWAiRQAcJDC1j6Y63SQYv9
YnSJqR8f/wwcsjV6G8YNFHMD31qEs3TQ7IwsCbFm2WltPLGYDzvF/yGRR9NVBRj3qXfI7in4rOcu
XfOoFNFaWCz2aH25TYtBjFoTpw3cQ5g9Zq59D5M71jLUjWDTQ4X7TO+oOV3DXTDDGRrX8SO3OR8p
PuSFuLQcoQ39fW2nGlELqtE08s1fdztIe+9/2EF4/Qjat9Zrt4hqTy8ISm2ChTfYH7DFyNriRkj4
vvU9/xiRuvZiObSi6yBGudbLhg/hHpkZ6cLbxUIJ6ea92JIyV2+RH/qXSNA1wc31vp5Zy1XAXi3R
7uPzonm88bpgxDlWKgA4WePEyJZ5YpVZu4z3eF5keVy+94TPjoeV44JlUxXsaaM12vucc5sZfCTi
mgfKdQ9LHTqfgkasXXYbENyqxo3CJgRoOu6KbBtOEOu87ZQNhY3wVKdFNuT6Pj13jbzVoR8OgP5i
h7EMxa1sdo/NQBVai3k3r1zCBPeDhQf2rL/HHuRO6UTmknDnmGu7/OS1IyeC+EHJKBtnP8j50GWR
mbWkwquSa7fsrIDm0+q9nRiWJyJ7zbL6otUXgK3y57cShgWWVj20FQNW7eLdgJpCV54/1dziR1f4
pbgKDAy8Wlu+m99QPZhjL4aijWq2EuBMmxHre672nllJucFmmdcy/BavDtFMBFb9FSclobdg6exX
DDH17/bMhHvIlgAblDl4Is0Z1O3kiQOyqPsvxn3pA/+3MfHUQ4PgJ6j2RgHrlI+UNoj/ZDAY6+I+
o8cfb6ZA+JnVzSQYmfM8c27ufJYq0Z4TOyMIq9UmLGEk6KhvwtXnelePfS3h14wZBCsLODQNN2mK
l9Sy3ccXYtq5b7RcSfWhWnv51+dMp7KuCaB/YJCnhx/qVpaX2Kzd9AApwwaGpC2l3A6pQCGNCJ3L
FZLE/rjaxcnWlJlS87/NsOziwJ3Z2BGBSPB8nr5EvuvoxenOmZHD2tNDi2FBdlhGJazrk2IrPWmU
Iv1yNWpadIF9Wi6OX4sqmCEnxmUSf6iOw7nnjZ8aSyxAvKUhsfCP4U8HX0d3iaSDj0gTXy55ocPX
HqPNR8tZhGvn7AxsHI2DbDBIJLxl/8kh7hlJlNM1apo/64NHnso+48sdKEKnD6+OmSTslFK+vM8o
hCq5kfrv+55YLr8xL29B6x27dkvVefnp0yhF4mYribpYTx5EOrSV2fmP+u3vs8sItu5LZqs0R6X0
Qd5XY/Bz75zfWKx9ZxSPYP2rgJu6MdV8jPlhWOnKPjOTkZxNH3hX4vgQipLyu9l3voxWo4QY/hDh
DcBaQr6fDb5UmddhyrwqKxR7nhFViLKiuABk47G09gIt5THcLfdZ96+zjGaNSbLpxl+QZ6Q4qhNP
iK/ciLRiWFcFcxJUjcfHcwaSDpbdzRQAblUwLDybILrYg+o1z705CGMyOGaeSW8euxTnTV8Fl/KZ
MRdTnfzIJvHalsNM81kwhnqLblsJT3/zVjXSuGHXasw5sB/wAzbEHMNudSnbbu/kYzDQPClcONS/
blNzz6l/MKBvRdlYHC5M7AHE7wk38HfxjEwadhrIqc+xNAPHEE7ocvbfVYbtsKUE57/5brCeLO0T
M85SOLUijrca8ORE6RX8oTyJFPi7owY9quy4Nn6TkCQ9vJgJHZsam9ptbXZlt1jjoEb37vG3Mewu
qNUTZiqJXmiDt9QSDAgMT8rNLPHZp8TrFx6BJz7quyJRNSX1u6Q+OkTf579RYvo6rZxW99WrkAZ7
tXdzHyOZ3/QBSAgzZjAAppXV7jFhyhP8ILOzX4jN5MkHVlROv9SD87RVBGoohzaR6kYeYbzZoVDU
ahDfrRuENKhX/cV3JhtEfRuvzsNP/5XpNdvO8dO9V+djyrYxfGEQcYvmsH7L7P8JkCX91A6wDlNo
oZrGaEzZRRugT4HKB3sX3n+MlWXhxeStUq3gDi3kUr7XsAjgeXp/7L407tsO/Sv+pptJv0drfLD2
FzQf6Nmf7BNQpEYYwavwOkrKXBTlbC5ffYbrbvkQLyFfwMo3noNwtm3vc5bpc/GTWI+9afA5R4tk
aE/uNO7Jg8yo9DPFOsRvL47igI8EjBxtO5wzOYifB1fpHDI8FX7jAfUTJDc5gdFz6j1qrJQ+wEt8
pq6VFxNhFll5ZnXZlU16WIYk+PyMSBcdavJpmx7nASsEaecLHe4FnA2DppEk0c8MhkMGAYskXVob
NcCycwL4Y8gT5v55DE5BMEfgP/jIhEkXQj9elpLf2sdsXUHsBvIVLUtHv3tg+EfBEpRFvXdJgH9C
5KnlztIbiJQPe3s5dAJEIkkhvLYxUqZ7rHMpnJ5Jxz2so8rRwq9kn4I2W+Rl9TGYjDUGfR8OypZp
ijWxo0sU8Kh1QKcvhI2tDxjOdPpJ/tO1FrJLv+2dbEBpFmbkpjoW/FNI4XUWbi2UZvZKBSgYldgM
9kz12pBweOW98pNvB0zFC1KzDWA9dok2KkByZXSdu2B4aevSzv55DY6d+j3FA1/jvcy4p3Tgp/J6
qAmTATZF9V6yCJh3mqfaddfAsBHqoztLXQkaMPT8f9vkM5iuANPGKSSkkASQysdBE5z6aruamhq7
qVsCo9+SsA5UYNjiArotQzebBURmTPF30/MfQFtLx4oFYSX2gWiyLTNK/3NjNnqBIwnH5VWHpAIk
2WwV82Rs+8/gLqJARLa1rCPhRmWsxR7uQ1VDXAUkj4MSQ6sTpm9MsQ8qBJWjj893ZgvcRfOVdd5e
7SO2MmnVC7F6QyzAwwvmchbEK+p/86pvMKZfRvQpOVv/dx5x8oJejTG6bI1gTLKtVbT8wNOM13Jx
RoZtv6pIUwdioRwUVF+3o6Rnd+tu6XVdP/m/8QzaH0rLVTdHEzDxlx7XDuws6NGJZAGudMub5YZH
eUWlnIaaj6tGFt1r/OaCt1PXB/Uy+Uz1T1dBNRpu1ju9rUelHr/zbWYydLo7PLlTN0jLX6jqzwJV
t04+ME8vY1FBhV0UBls4IG7n6nbV9ZZUyJAKn/AQ/woA9Wyj8hQHYam+JP8z6xQnUcSA6XvfReBY
qmhwnBxLB5gJkYRZ0KgO/72v4fnAjwyFggE2iUVtyrpuvn4FWzdy/9k8c/8M4H+3MWQtfZoHIIjB
S2IOcMvSPQMsHiHMccVQNF12+QiC+Tffg+TBzJs7CTjEt7ZWn5UCsw9oU1kU4O7C5sch18Z0rzhv
wVu356JJX7HCYF7WlNlXOKR1q/fBWkGSvvonhXCNaqHKxtHvVXwF1ojKgvLm44ud5XsHGkiTblfS
U3UacOU9mDJUbwwhr5/z8vB/rr4qscAKC+yNWDu8MEVhIPE8P4PhtDDjpiWsVPAkwKix6DYCENF2
TjezmJ1gZj/X2VBzTvyWcRtXGb+UHYo07sLIGiDLLEqQ8kQMFeQoVtFX/08WBu1LdK0vgXhEsvGo
SUTs/85RHNztkCzZTdGtOxXV9L2eL7Hdn7R4Snj/PxEiSmbhe7n4vPHlhG1TdLuBh84iDmt9HghP
u9mq6CG9Uo6XFX7q2+GZpjdcxNm7a/Vw8gS9VMpw5PWFGRspGzfbb2cHge6b2xd1fP4278gY6/7d
H8lzmglpc/c4oreeQQxttGcibqFEx4znwTxAIz9Fnu3wqwzz1ctdNhOQdHk7opNL9IKAIP215Cr7
HzLMj9X6m3kkyZD1cHhsC+iDf3cadgAYiXQi5eHYZ8gPqcOwRqV9j7q5396TpD8Ny5TqBkDssfPk
exHxl/Jl6UoiNNF5VS+uQGVqlhV09wVBH2yGPBeYB650HhOicAaagprc8a/qqMbQieV0MK5XpdUT
rnQ0kV3MOlsioXwTNcCrFYVY4Ng8ipH0bqKt2SGRdCbGpnURj7ZCLK2N5neXr0goMo7/qSYsLn0W
7YaBNIGMlFePv0mPJCJNZ3gWaimn7PrNn04YYQu2rnpAEgdgQy4KWk9oOycoDzDkqc7WgWLJKkrx
XOiO4+M5EjzqmZbZM2cCL9XINTnFBi5knw1kvzmXwWrnZW9/8y+EnUh9RlDl6RxtCIwMEOKTY4jT
JBuWPQBjULvx1EiOK/SRGcweg3KHSHydYEg3Jfm1/pYTQrqYtGrUIVVb9LDwcZA71cYR3gTKi+9b
AjHcB4gk56qsiInhCUhIkgbgGOYZq/t1v09BTf+fkDB/7gymYbek/lrOWF26uZgo8Tm9Qx5k/ij3
NP582v+jOuawIEaTp9TsUXahh8m2qxi52a9b7OpbQgFYHl86X3M3KNAmGRjxUKuSAaZ1jBbkMuGW
16faxO0RKViPJDa0b5+DnGaZm/nba60CUlxF68BwhdYZOkF5EXuOqERFw6SMB2R2lUB+yGcaXihs
KNv2vbejzGviNFxHwDsdOj8gvPbWrZngVcACz6Z9zZyu6ccnrc5VRvlFedkiN8FFPARCqXhsrw0b
UfzhrRM4WMdC7/E6NxP4crewg8EfKr/NYwtClnrJLi2qxO3++3UqzNiHsy+J4VNSz1oN1uYs0qeZ
JT4B8GNZxOVVBxyzsOal5no5sJuC9dKZN9PeP194rRUhBURDhGNYLxjjknej4GWMuKuCqQ+R0u9E
xENaq5Z94RXB2Pro7+DQvuvWdd9C2uIyHHyJreucxOYUu+IfFOSwI9t/9thFFYjxmJHBPBuDfWt/
4R7tTF9KzOefgQnchn4vF5yFImC54QmowbU+WFyX0yeAeXWP/x/XKpSB7PxuE8gY4s74RZ9CCMni
tVirC3YdxjJwyiiP1rL2OJV1YhL6usz/1fItkutyLXOoEdET/TmWmvFv3nHcvEx0mWkY9NCJHeDK
wMIG1vh0EQBROxNbJBweNSOTJCMwcnt63waKiJFbWVTs5pCbDee4BTzwV1k7wjdeSvEfRPW1RXtI
J7xhHtMoItiwrzRv3jEruqYjyU1BK9F7eFubA2KWUhzC21TU2ZvHGZUql4s+ZK8B6Te7KzGN9A5W
A2+WOdmcU2/jAO+fQ52/6dvPVzr8fJ7i+Bro3qx0ahwMPw+69IOka6gD1yfuUqFoGcB6VaA6nuqP
pwXujHTMZMPxOoVWPRjXQYsKO/JL+StVfeM6vYwjznctNwrS7qTV8+QY8jWg2hKlzBb96mdzd7GZ
b7b04Qvyu71QjXGktAsTmtAyfPk3jzL1WBknbP6wnMvXGaKQfPEIZK8m09bKNA+e9YgMM6WzfXg7
HWKtASnGmohnFtnAkdR2PxaI+RJ/lINZCa4YJTXtMe0dHVRYO70iYq4xL/w9ZROnm5EfDFgaPFD6
fXbWyAi7Z0n5Nc2kh2S/JGQjiQ9VvdLfbqPjAAFvUgr6HSFd4MwojjaGuOdNTYBR5Tua4b0J7G8G
VZb8w+3GfjUIIbguHstFaJ79yAYJFQMeOEZ5uaO8gv0H/Y6cj89k75SpeIoAggpRWmeoCWqMKJQa
4g+8qhHCCfnXiGYpR5Zja3FcsLgREPw22NgsFcujlkAsvVx/GJVBHGRZzE7keS67591PL82kpPIO
cVB85oJRbzFjB9RuacQqOerEMjxPFjZGGUqW0m2ibNfbptTQdTgoJtwNNEP7Ykhp6p1RRTe8zxj0
qrwkmj+lu8PIlD1k9oWErB7fHH+D+hTXx9JtZrFyl9qsFshmPyTQNBgyA9fWzhUH8urXqtn/NvxG
EheW+izZ2HU0CKVPtivWhcC53Qjf2jJdpx6GRWxMWYi+hHXn0GbAhmBLe4vdbDA8YVuUTgFQFX1W
TtfvpKb2y/NruF3XUh5YXiVVZ7WnGhXWK8Cv3zFpIlY2lw/zpBDfjmDw2HKPrs/wxkkKE8U46sIc
RgprKejT0InutZEn+dOXDuCOmCTCVf61VSWt8GKyEQ+yUElVL6duVqqWtjdNpiPI56QmSrOtneti
l5UQr6blaZokrFLz15iJcl/M6eNvLaCPMvZ50URpvRU3/ez4SuZ8pIhLffYYBcAEpUkoaZrHuRla
lsmpvjqEUKAf+tt/X8ICcy7Vbbwsz9U+O5pPFvHUOTRgQVaKeowTBKw0FVfPMaBC6LlB1ntOzl0+
Tyq5mrh40L59s/bj7p9Wdqdrf50UGZyzGnBqeo8ZxNXgFlnqZcC4g35XgxdYXZWbsA62mDgbZDjo
Y/+6PzyTeX575MAyBQK6tGz/STcjybcm/udorRHCyc8i5wRoYJk8Hx6qCahIPZ2GiSKzQM0UOav6
TgL3yacOHVjgjE/k7snRkYa6MUzux9yN6W8t/Okx//7bNAurCIh1vV/9Cvc+i1GFOdzaMkIZNjIj
/SvaITgQK1JIP+Vl+XLCWz8EzeivCUxI9pVqakwk4aGD+zTV2uk6BWdMet3Udwf+nZYIlewNmK1l
amt3moI7vayBzJRJVOqiiHgCg4DJlhewmiI7L9wXqa9LpSdZo9V9dWSYk2KBP+2jQCx3JL3EfxnE
40+Xn3p5Q2zdO4H8+uVGq+bq8D5ULCB79IId2Ni7K4bWNsLc+TGyBsAbXt+S/0cIhu6lGrp4Awyu
8elXmkeqf0vcd9Q1uUd33BvherJIEjWqypYiDRRTsdr/lY61W1cLxFEuD9mv/repcPEipIvz9s4i
8K0QltUFOeTJVrZx1tNzH+rpMUlOhSqYCWcKMnQKtAIZjhzu1I+KxnCUSNo9KAXWuYf/g0xVW0G/
Rjn2ywSMgmg0BqorHCtV1/EoTjV+ihWNpz+eV4K6SPGqBtaCQ757soGU6sG6cShRULdNjv7u5CN2
zehXYS/RbyQrPhlF+Kqp37mghm2obphPruDDZ0+1xCnkvfCK2DklTdWQb4EJ5/M8IUK/W61hX6Mj
7HxYAZ9noj3Ub6IY4kPjEL3vRCRduKcTib8VFQIl5TfI2mCmfD/gIdJPgsBH/+415DdQgvjmgqt3
QCsI1539MasXtXfeJolnqMXZPJUd4hDuvqhhSSpYDN2R8uLzcJcxAO2R5CWrnP2YuBK1u4kPRbcL
MKrQ6V70Ibhm95j0aj+wlvqs+xPqd4JlAoC0QM1t+qkCZ8rmZHDvm9DU7Wk8QyBbCWIMxEeK3cuK
vKta91dgYN/1s812pSjV+nxAQGxeXKC++5zp4Nx77RVISOmTr9WzquCakPR1UB18rkQXaRHFb6HM
wWvXbwF8ew/KXhuGpc3GuGUl/bZDVlImxtb7BE0AL9X6cT8G4mMugGCWvxtP2+NjitLQka94xMkh
nmY1Zuis0NiD5kTE1aNI+aHO1ZV7G7ychb0PNR5enn64a3TEKkNAroEOxcjQirVO2heEVlCMjios
KGSkwLrmx7KmsKGxbird1ruD4vYfopoBQwBh1B4VFfkEEl9YHgZIJDVnOiNoKNUnf9QYnrplyNA0
uwVSfC7bZToV9UTjIOSdf4OsgXS7qNimq3qZZ/ysZ8dyrJCY3x9NcmHVhdT1gnOwk5nHruVS08K1
MCpZ7HEor/FCr+CXg/chX8JZ6DmD7TEonNjSv7yU00MvDqNkhp++ZJIXUOLOSAeh7yKKx/iI7g63
fasQqFfXwrT8VBknAEfuQ6QrU/tlEdmf3nlfxtKJ2UpN3r2x4bHoPirfNquwxr4UejO7+r9vebxV
F8UFexTRnCQwyYFh3asAwKubSsDKUEsW/6q5BBAr/NbsuC3JRX/iUBxUT/5oz2mQI4bEKSVdHxlC
ERWtzQmrh5Phs9j7G7TWY68x4kmyyVOHQb4yZXvU//2V9Ytz3aQ2nLl/1YgFEHoc9bu14MVOaEaB
7dIg6nU08q4GvFgCIfxDSJzoQPtQyT/kxn4c+qQw8024kkRmXs+CuFYTIxBdA8gpuriejPpM7NZw
5sP2ymp2LfDtPOQhGugq0m/7dH1qWx2Tfw67wCn1X6oLVA+z3K0P9edkETKim6FUAUr25Ax+mi6g
GRzXJxnltcTfIrQOsfKPjldAgsw0eU55sovCLDgwZta2c2z6IU1Guis1qHlfaydq+w/vJFclSGhl
ZUDD3h80U23dud6S5CWATSNhkRksr+0Ew4i+tLXUQU2u6+6e7MkNJDHgTQ7o7MmXfuT/z4OocWcW
lc25lvnBnoNTOGmxKibYGDgDtDuej5WfLcMgM6lBktgQHOV8QbP4B06PuOGzeWy8sgAymNYzs7+X
KVVR6MiVTp2P+01rzBlVwbUN9HgjvqzL3VTMTZHRtcx4uTDj4nqNVv1k5CkqgdXi1dmuUO6OK5Nh
sxx3tmWVzog4ZT+2/8mSK3ytMsR13to92QNdRgTbeXSZ5yYpeE2ebY70wlKWBEotrzw4De1eUSbJ
60/SDqPbqYegaOaWjTCK/gNDY+dzauAEkC+nTouXGycLPSWDLns+3t2En80PNc/K+l5fzhyVWsZK
O+lPRlRtdIwa7wPJv0MDrTj6CiNP/aO7kZpfMqywx0BdxkUBnJ2JlTy23lX6zTNyjop8bGOvH5Mj
qiUIrgdvcbjtbToUz72Km4MRhdPP96K+yySOZj6mPz1Deh//TrIPl1+l9B/Vw20g7Tgl2YWih4Tx
mSLTcK3bG3AbqH3B2HofwnxCKiz8U7V4aORbEBJQaXneKIIbcO07UahJsl5pVtTbmtEnbXGkWOEk
w/XkfBM4hmVEx8kwiqJIktP+t171eTgtWKboVkI/YmM4+BkTKGfSjCpSNfOh2Fb77cFK3QfYIEy6
tFym3h9Ybg4N3Eq+2Sl9z8RVEB0f1B1xXqFIkuI3wIwUym8Dnkji43Wa8CYYRksaHX3nee/n3nH1
+tuNnWHaO6ItoPM2rOyjehIzboPC736W4pNozr+aIiZjRoOPh/jSWjj1QVOmg+eDHpH6bepbYTAB
SmHpGIjQhJieZRH9spF02wSwflnFqLDoPnaraYJ7k4kw2cSGLaXOZ1CXYSFpXPDDVTfmwXakRGLY
uKMKt+Ja53aTx4ZvAu7CfALnFUPmCJyJftLA054/lEUCy4cgaTfkwmmXGqO5U0VOM1bym0L/mtut
4y9HGgrI/r8SX8AAwpkPxrcfEkt8CNDJiXkAZWqiLxV22ACs8q4YuniVLizuS/YeWT92zF3D7n/k
4NbnOOOYNAUpwERg8TNyvjSY83KItDclWF5JfEm++bAaMPoVZCgs43BnaEjGS1mUMdVecYmeSLBq
6OPetCfokRgPePxPcXfLgjvJcOWEJGSFtfHmqgGUln8fgSfJnoGWqmTU4Wi34XpIM1lwr/6LIqQd
cV8v6McTemJxF+aOhz/Rwc4IvMsl6gIH7ulPVPGmiozWKoWv0EmJn326LXAjfrpgZy7JlPS3lyFZ
iPRmnQ8S/el7rQB73j7+ZXrEeE/fTuBKBb/H+ShieY7LxCVwcDFqUQhAokSapMugnRgxhRPpetp+
wL7m9DJkfICnocIyje6t15vSUancrab3PDscxBX3HCl7LiA7HF7Uda+smdcrNzxrekiM3b3BEw3E
uymh3lSbdwW8SRbz6qccTMYv3RCazXMUqahyYFU1NxUuVgKEdd40B+l2JBmK8Ul1YySAGQSs5T8D
afFQOL/tsdn90ySTpr7O+Z6tw9jAJMWhrwe/lgpUlRfZN7xzXvHGhYZ5Z+Ei45kMENy0I+bmC7jj
6vq5ono7SFjYnfJ62fruw1wLZmFPp0CjaEqU6i6fROdtma8I6BMxwVE4HDUs4S4xnZHTbii20I4k
uyGVtJyKnT7GxSMXg4m8QBh4hpt1/APAMFtLL58rsOil5L8/0YCsil/i2EwmqJfINW8I9wap6vRY
JkjA3/3gfducfHOY1mE3vkA92BMNwRzu63omAnNgdW/PXaMT4mj10MOBTHhJ9Lp1RM8uaWJ7L8zy
+PRGANbGdls6DUqnRJ6bpA8Jyf5Ed8xmVfXeMoaE8nz0f1MNRB/eZvD7H/oXOof51fZcUE+Vphnj
Wal7250TQCyCwvSEEgmdOwB8+gqYWcXU2SCqjl7Dtikrctnc0rsR+kf+/D0I/odOc8goOeoi1p3F
xSvo2w/YJFOxxKoI23g8V3WHkWdNPDAg3RArt2iGp4d2k2JaJpDAyDhSZ2s/aKdZdgCH8h+/9tfy
QL2pJYovw7aL+JnRIK8+jioDNPdVym9YwOHPZtBWj2TQKSxRAOVqzoOHctkuMWHc3DKTy5kbX+R9
s+DSjHMB3fK6FfBaCtixIB2uyrf+xaMSUctdbzw3Z49zWJPCCPRPwLq0M4DjIX2CNgv51AmUSQg0
NQ4QC4B6jgekMaw/F0ueP3ZGxALo8E70GbQbpfi2+Vi4Z8EUTvep5aJ5yj7QBqz2A51PG/wVlx6L
q/3Skd+yibZjzRNJm+8yikJP+Qt1uNi7uyImuy/U7THZb6bcEH9VkXrhutnw4rlK7bSmTK3vzAL8
R74nac7zifONfBF06X10d6gFbW/QlIu350PLmHhParf2xodfT/rPnIhsaKq1rNqtv/3TDfROt7bt
0popIbsLOpYDY5KQuZ3JCthZpifShAWfqCCXPkJ+qBX6F5yKTVlZqRIfnutP7aLGl1Vs/AUpGeS9
vmrPETsuTXrwgnLXmPl4Ftenp0/0vCY5rkT8QWo6LcqAyBUH6JUDQkOk298H750SUdfJXx8o2Wms
gNnZSkf69mT+H5lOhzZhD5AI2v28kxjH+sUn1RCrp0Eaz/3Byk4r0Vg4SMJnYYSVlA3uqtAkb8Ul
Is6acw0JC8jmPl39Vy6DkrQ3mBPQW1qHhtnV1OJjtakV19BDc6EjqYtwSzTnDJ9NUaKRgT6jCaM/
HhuF4DCZzpgIwg/hzzmK0sHv/2dU7s6Oz7v/OsDzPQKBVqcwBVSzOh6J7ikGexOgMfeaFOk6hkbW
PWcePu+y3soGEiiOZ+Tg2IN2/k0EfWod4lo8zYkfIRvxRceHuIbRnTCCP7mK4OsUYw+WUWnc1Fpc
Nnisz5VHnuRolXHqpRz2jPwoyLIY0ZNazuNnqz8vljZzG6Bl7kiV3JfyfhGD3QsRAGw2lpIZ2wDF
R5fuqHqveeEH29MQapSNtS17i/VRd2H2CHJCvMKghaBc0pWPYYDjLzlN3A1H6KbpJ9/pODlwenR1
EcjbY5WSqOqMlubmxe5biFi+XNCNdDpaEGSE6l1OrV7qEr1hlaNCnF39B6yM/uYTR+i30Vl7TnMl
qJRUSrwpd0nbi1X8bGeNdOtr7Yam04ruY+c975EkRP+CA5yCLqW92dieEr7raFM6scyfrezEGHlw
CBO7/9l8Pr8uzO6LWRAPpXr5TKHiWKvBUsj9PILYMAemlzgB9lRpm7tpD5bSrrDOBi8g7JLlhLVD
mxdpZ0WKTxHr/HxhRWvtI74iFzAuiNm+p2Jl66KQxxB9sHJ5x72JLaWelwLBI0SXbuf3QouGeDLf
ZVpbvZX0xuyxSoM1JB7do7KstGsXAnFRuRnUuuhtM+izSfoRtJB+T83W6BuzRJm0Io2PN8ijXkRM
uCmB0FilVpTkkTZGhyU2+aNaiVXop2SpZhnTg1vGmz+Mo6k+kCoFJKZ5VYHRjupnBHfx+LoWVcM3
gGgfhaB88kyEsc6elBadVfyBN+wEFUPStr6rPUjHzwk35MWioBm0ZjkFpvvJ+MkBmkFeC9Dp5gjg
MkYbaKme8JRHE4x6T4S2RmK70D73/wZQTU4DcSaRtDefo5Z35J0p75jRm+XzzEIEtTHlOvxtAPVp
phhSD1TtyzFYfzhOl29HlS3d8JleQhGKMPaUA1P4vMsPoLkdLnUzwqQwcRle9zPB6EX1WHDaJGJt
9bcly7PmKW5juyea2ZA8Dncc0zAIZ8cieaJ1JOp8VzvV9Mno+bfbgo3GGoLmvAiugyE7malKW7Do
5MU7j2HJ99CNkZo85rscUiBkopPaRjN5raTJzr4ifWeC5DDT6oXPkOK6CPII3XUEvp68bxHPSmq6
POMXtCs906BR5tezg4Z0Dvc5h5qK0qrJPJTRm3Zch1rWsAIdf0OGq6BwxoSmJvcntwN7wnQQmJVC
R1YNnHN6de2uqRksz47zk8W9GQCu0CUx81XmJAm10pPx503p/8rdLduIkeg9sUn8FkAWvZttDhWd
vym07ERAlCQNrZjGXXDIED6iAwEiWNrkfimcQTjyAixEcpskjZ4eFKWtAmVy1JRKcD20xANxhimJ
pBjRZ8bE5+k4/+yh6499fORMiNBSxOV/kUu8VsZZE5SRVttI7aR2GzMHIfIoOfsjbpzI+p/yRO7l
OgF505GxyyI9w2NE0mxlFUk1Z2yaaOzJLl072oihan3zOm++pxU3x4GRuqMG4NreSmsQMBK9mlPS
O5cdsVeyiSG1tdcsW0gjvzpcRWxKcklbwmUxtDrZN4MA2ni3e1No5TDd3oPdrApQrk1Nnm6L4pIm
H9kIvoHMCSgqL5mOE4ERRzmoduYxSz4JL5e+21arVUR1kW19fiz9ZBU/5OIkZy50KN8KeK6XxEri
zW+sY5s+1V/h8bhM33r5X6ynnTS9DeVRl7vLn8I5OG/TkAoGArR6mwMKMt5ThK8fh8TYboPTjRq+
RV0IDn9Q3faKnQ3v65WbHObdLnJB42hdWhdCEcOzeNR/nqYjY0QR/RcDNt3tdLhYlIEaZRDvmNzR
ozBD/nN0wJvOtsW/0OnusQQYzg+Ba6spsF1e2s8r8wrBUJBsnz7Vyu3f2WmV2ty+wNDTDxf2BMMC
TuxAsRiU/52nUcoPQaexpwgwVrnoyumvivzCA2/thbcDzhOz2iJMbFehvL5N//6EPzF22OaQMrDq
8g/Z3IY07GJMGTGyfgh3u6bUL/lDAuctK1qYHxLFv87/Y3v+l6wASxZPcU3RihUAUxbJ2spxDf6m
NknpGiTICKaDU1bJpqJvi7xEseBBbPHik8gxX9Prk7IR3QwYx+d0HBvUljKpixPBLFF6EnELRhz5
8jkVYf66XQdicBkauPE6dAD1CVxWsDpkYMtU2QEil2gV6QbDqcgWijPj7Co0UlzfaYi8gqoG0HWq
LGySaUvNB4nwYZX244Yg8sOQfHIjhK1sWO7mlJo8h3hVQcGScXMuHvbwOdLgz+AsJTtKDXe9SNr3
TrdNIQaqU+XTrY3s8xdr1OtF+wzueiof3SWAjV6BR8frcR3I7e9dm6jww6wrKmlWVPeisB/eou56
tRvXkMC5lEB3ti1NatxmXrbXq68C4/qol+e+TJqvXXpSFmjDUmzXjzV4c1ckxGrtcwBp5ZslcJow
6WxaRWj2fgdgwkuwzmdsm9NxS+h8SM32LXEItfU16C9sCuzHkJI2ibNWEt7wfd7NIvA5z1e3yhxi
OAqcv/0La+i4yDAWcNBMiDpLx6TYV8Q2JsTZrKeeehjU/A5iCRyDCYPddWEM0He8mbDR6MRZXsFC
XfgXcIXqFKhgP1iPZQ2ATJ1OfTNojJQyUaclv+MaEYTLCb9hKrqy8Mhls08Oz3NibkKPtSpHFYT9
n+K6yTLVEUOn6URwiGmn+FZYJh3uO8xNr4b0W4q2mctlV734qy2lE5uI9bMDaDfBthKe95U4k/9m
gYxSR5Se6CAGlSNLfxDBtScVSDjIjdWdAP9P7BcKwb48J2/rPfdBdutRkRY3s48lcXymaFdpYzyg
TvZMSk8pJWIsBBmz8VkUeGgrTCY78T0rP2KB6itqMTNMSeK3aP4+CoQ/AFZshkaCtKGVRG2t1QZO
9/VDsIEvtO/WO/snQ/XjcQp+iBU3vNVNpFVivz63BHVef3F9p5ryhNEwKl9zOFN8NMDNdiqleGQv
OhILALhjEHAcuvOysexLjmhtcPpju4tZh5udLDhZPmQ/N+bvx/83niDR3NjYSSar4Cfl9hCZn77q
W5zt6fOEQ6tgmSCUh+AwWmmO35YS7nAWicQVf88Bd8WRO4PIueOHQ6t2uVL28jABL62yUcT4zGwc
/vFtAFmNWCb2Mbm1CmNsMHHDcHc1+bC+/nBP55rGvzNM6HOz4kPwyoiXHvUYJZPI50c3IxD2KSs4
b2kgkhEoaI2e7AQcWX7XKdavcPeUJN22tJz6RYACR5kBqydcZXIw7qi8RfxXVGKJrhz346NkZ9s8
8ztukEebkJXEnUoQuQTWWu5/B7g8VoulvhsdMN9ahtBXCGOnux3I37E19NLpkzxFGFJk0L1iLd0k
H2NIY20NsJPja7Hiv9QergjbYUgNKXGM1oITNDFG3+GOVKFxllH/BMCRXuI4FWaQOj4lgvIsFbUL
LrSdBIOut5Pm1SKLsZ7MGVTOu6i6fHjLzsc7wD6+qIjQUFLnnqhqrKjGmmy+YtSmKI2h+CRT+/Gn
iMAuHHSv5rVV9/XsGk1IjP9e0l3SmcozDzlWsVfuAD0/vf81cu6igNfqXiLBpHZMIES7UgqVQK0y
E9WdQBBZw2SWvBsqkn578nrl7kf3RqT0j+E+mrfQ+xvf00aEQPor7gHaZVgU1Hacxgp+urWIYpzU
76ZbakMr4nQhJTBUy1c2QQMLnb1a5Re5WhAR+eUPKjueEBpfy2jrcC4Aygp6LZXqBqEsR4yPJ6Km
XVptjEm+6yziPAuXVo6OfdzFGCjOD9yqb/c3Q050CEjNsajzgEXO7XEwgI2+DTIMpC+lhxRdGFGo
At5wUYST7Z5osZ/ATQ8ZzXT+7EOgTBpldc4ACVmSjIyYNOzhHE8Ijad1kswnHAPI8AWu3RxsS1z7
qEQO5X13SKIJASSt7bgJNCBkQGOJ5hrTeY+iNj0bXjADLkASZMr8ijNwVaPW4rejxEfreCHzGrx6
dgeYRmn7yoBPZ7EkLedJkV9I0aESPflDY024o7Oue5kTCQ+wczhSDo5I08FerJ1CZsl2dwBVTX7c
5UnSCgOx9Su66Dr/5rIBo66A+qXMDpON1wVqg7SLZ9GUrQbs+xl3ySPKlCjprl8D9JVwRa2qEsI0
pomVXJDu8G/kWlHVmybtmCuHEXSo+3/tz47TpKP+bZNnXi7f88DhJcqcZZUpUydr6ZXT78GMPjdU
vExeuSQTFeQ3wq10PoctjT2LVDib6eUshcKvsQgXk09yk/3UXomgDUyILWBpPvcwPfpNjQZQBiQ5
gvbhPtLBgV8n3HVlnuAWucse4oSxsgM6IlLjHps1DXkIRuvbbr4+aISzpin0CX3b5ZT8MUjXS2y8
9f2GZRCvPMFjvj8aye2eeYkYDfU932krSkvtOL1T1CoFavj6fb5mpCRxVNK5B99uluPitP7MJZ9M
xf9pzW/eEo8Wxy50kV0xon7gM+/eTIB0XZ7+VGpF2e5/ytZmiRPLcN9QyCEBsvqlZg1MCp3Wi0Yf
tv1VwC/PPfz6yaWOtD1LrQL/aEj+TQ2B/yd6999cePpSjhRUYwNuJZEjDRT1TuzRyBR+K6djlXQy
E+29BSu/C5ejml4HT1i+zMhLV7nf7MKa4nzY14VpNspbDTCyZTUm3Uwwl2LaRWlFxRqU3re+tOis
bm/5yog3ZiToKXjqnoOHEAfF+avoK1PhkpH+xt1cPEGSBElFlC5da6dVrY6M5iMRTWd90xJdX15P
sa41igT845ViiaPzFHzSWEjQs1Md2rvGc4Dk4npR6DDd10i8XvM3NuLjo9wyh0IDgBD7VHnAoh01
ZdJeSHLJTUD1UIftH1V6BaaTZY3GTF6shdGUmBWTetgTWQ1UZwO5jSWJdIQYgBHqS1t6UPHdupRI
7MfTFSXE2FNuQxAGOIatwCyW0PbexGQ2dPBTp3q/6bXmv9mFyl5TT4THCIYFFPO7rlGOGtNvMS4n
bFpYeISdeQb9uj+K6vKmZXsrUPqSKrMaPyUyHnbAL+8+Z0unjkNKqdMomOqsOe4aiGrfUk4UkmFM
6qS88UucEYTbZLAtCQXeCNz+lUBtxlxRuUyZj8hgL1+I6j/EEcQiuzqRIpINL6t/bjwBSYck/C0T
JR48DR+N6zAgyrJnYjK9nOIM3rqTN3n4H/r3cqX8NDL5ub33iXIPVUH8lXgul48gcysq9A9R3fBr
QNy6echQR9lfQeMQhmjToz+THpLueH20u8dXvKLmtrkfscnMJ9E4O06OMClyPJehDZCm8ueGcEIB
V7n8yyiD3K4HqRjFAWF6jGkvy7UveQ+WchmeCty3P8f65sgnMZNw4CyBsF1aAF6K5TId6avnK+gG
CvrtVANn+dHd5hFv4g1HcM+y7Kq2C0R3u8TOFn00C3p25CAH1EsRWxYyUmO9/lzt0vaMV+9691Qp
JZNEYug6LcAWmNw9dVb+v5iyneyJ78aoPEi3iK5dwLOSghKG8hTSnPCaUHDaxHSwnN2iCh4Oyf9g
uEzWZDQ/MQyjvtk3RLJrNSW/IW7R2yYJHje87ieK7vGnvPLPGQyZiSJ1ZghXqiZSntjec76ngTr6
i9kjxLp2OzpfFxFFyUFvET1UH3OyZfVj0bd/cJnRBRTpGF7uVUW292mrfUxQ4yOpEfMSZZ7ktXZJ
8MvwQVifCknq5NzJiVPvIfZpacG5FBUxv8UGnXtTgiXYYVP1Rrdcg41Y9FngbsJwgYlHMJowGRMb
jZ8QuajqZNVRYzggaxRE2nDNCbs5zzwbyihTYruZGKYt3kqE9eXZMYBRM1TGvsc7J8CWmeoJoRss
ibz972VBLnWsopmUEFo1GrJ4oXFH6Yg6DWkPbgfH00tt/Jx/b6i4aXoRu0zvn9TvBCIY8qj0C1Pp
UcI8o7BoTBnsCYGNbClaEY0oAj8Dnox8Tqm82IOFQZLQnT+oJSV46PwqTYduVPseZzqBes4mKVnQ
bzyD0c3JVFsTMAsOaxGc/7ICHaJEnAxVD79m/sWDItUiYeK2judnBWH2dkK5m3scyU3P5ZJoOZ8y
OpHm8Ihb5lMS4zdiINCGJj9zhbYpHJcXJU4I4eW43Oqe9XjfyKwCqRWdmpeYqGzQG67FWKR7zOG+
wDpbH/F+QIfCOIJjqH1R4jc5opPmExs9jkJ4ARf0ZBwIwOaemz32dZTJsz0m6/t8r1ecXzao9lMk
A8BoDf90ixHwKtaY92m1e8s0l2fjfQbxyttUITucK1sT12J5jCOJtr6TVU8pB1gkumrLLtvAh84+
ufO5LRebuEUEZDoMuwaGnZ+ztmcv3wGxVB31XGJ5Gw7T9ts2Wnojt6k0Sw1m2xUW7gQnHH05g4RA
T8fkPdTojOyhD9ZwuvQDqKiOo5JPRx1JlmJo6RJmYcA8k2pojm86vQbEsSrRmumeuBslK7QRD3FU
nYGOJpAFa1jaqttGXkQOtHTU26V5mVW7/a62fUDCV5Ei0sUcNHgIxLFbGYhuvy+Xj3WKhwJA13wg
7ZPPe1PPjIMO06xKNZUY5hi38KlypdMIWYIvM8/UPpkPs3XIzPAU58iJBG+FiVnc2A4ecQida3In
FAHipnM0J+for1TmduNqfbbKjP0lbtvXl6D+MGEt/3IGzz1FaxUQOiNh3TMnCX+cQq+aNlMmM/ys
wkWfZ/z6uldJ/R63Ucq/IhexFvElc1sEVaY7pTx4ELuF8kppLLCnr2KOACBciQDREIDG0eSxrSmc
Fy68U+ZKlRLwiwvG+id1Lh6re3JOaThjvEZnrj7wSLEiS30mzO3qywnuFkHTOrQeN2kwUvQCdhfS
Gatdez77fUPbXiV7UwYYSwxH/scEpKdSOpQOn6gSRj+u958SVP9mDcHI8amqkL8qD0N3Q2ttIA2k
+vmPORj8pqCN6xWG0wQ0QS5womBnqS2W8R001vDWA/GgqQOlSRdrcz+m4/4r2pIuEbocKjfT4A6R
19M1Qx52D2Gm0rYWVJyPLTUHTTskA1w2ryE9TtsgZa9Ah512F+prI5hr/OraktRDvXNT9738yTDp
i5oFblGOeS5Ss9coy+QaxUiR/15UMMph+WP/X1dOaRAxVib5lrTU8XvkXGwJZlt87B/iplrRjRIS
vsA9vdI2mwG4pJXLCX7PWeBdI1vzzPQ5Yx3Tjvi+uPgVDwfRqWZ6Lkj9/tjfVdJjrav6qGF4RNB8
pdrczmtwnimbU/ppMCC/JMY61SdIxYB/p/1vPZpNI8CyvHvgWtNjFnDQAdpyQW+FETHtPhqyY/aW
kVYVnXDWAtanO7YLap6QR08k1ituod7GyUxAszn7g0IikCVn607HnujMQKl9O6qLHfPGOzJrORbg
CIHJ3DTJgdG7fD3P3jx8i5s/8Dp81sOHxXDhluObLP4UkuIW68BAW4J/bZeh7+bhKpF2n8mVPd24
eisDgMpDgYfcsxYp/0PiS7ym6bIzzNTQOdxXkFFewspQEhOSL0hixRohSQWz2A5jmuOGlR4FBfot
HY4brna7FsMjq9eMBEwBEd+mscil1UN0Mo5LqPeGNpvIhHQGKb+zWKsu3euStI0rEd5a+7WAL+qY
A0b3UQgHyfjxtscSU8SSyTr7V41st8ZyUtoKBW63RUVSgu8dh8SzwdigBDsyr9rQYC4O3CUqOZMR
O7MAk4qAZ48MAtgGlXuERS21SfuerIegyxFplSvUtGwavEBBtRnyzfN5uHA3hsE3LC8quf+V9iON
WPsiyOVZFzDyIvac2FkJvbHM3ae15HRSukT344TOeNm1DhJB3FPRsdIoa2vQ3EoLD7hgExSeRxTm
8WvfyWfurefisQzwGYETkYKdzDGAJYstCuG6JBhJewZ89LH0nK2xcee1SZNnjiunYFVOfljighLu
tFQO43YBqhvUWrn96oO+ju1dvTZRhI6/H4QzXLehUadXkR5d0XAjAqrNJSsoCffjPgfeaUQFTGo+
9XTVGSHMeqg5Ro3Cm4Qd9p5p4a8/vg4Rlzduz7gHc4Pne52KDCjwlDHm7dI17P+rKB0bFImshD0T
Kyku80spIQxO/VtuuZqu9RqvPNDIyJ17VV6pIZHnyMF3kvWiXU9QDgErdUcoWypuGsp+DySF17xG
KqcmINTFrr+MvFpV2qFYj1Zhc8T1hu+TB5MYAMyU9Y4JK/0jk9xbGddfBVxBZKhgWJ9ca/rvudo8
rr1RUn4IKy0H8tg1TUWpXkEQl/wUkTEwqh30edXJUV+YEcd98ZI6z/er5NOKamcz1Nk2yxfM2oLB
OXqIUAqZbjRH5Q400px4VQZLeOixc87bRJbYWEka7fdsSQL2vlCRsNR1v4/0RZgQSr/Z2lka4mYr
upvDJjV1AGnQrcrdHpFUHw2fGQmFqxA2hDbT5CKmNakSdQTHaRIdLyYYK+WUgRI9H0wQaniKHKqx
0UbJqAnE8M7uDp3sGODq3TZfG5wiUQ/GRrTweT/+GQvZZOXqoVHuoVOpo/orEosCiyTs2QLN9CCg
d620/Hn6Q25SSLkQVszTdHesbIvx7+TYfP2idEAkqoSkwoLKkfJxpDFD3TD5sWzXDX2M0kY/JgAx
qx12nc0cgFudSbbBzjku/djkVhxgsHLIzbu98bxNW1ncFUqWx970zupqJiZLZfWVMf2NWYMN/QJM
G7iJXdoobAmTL4nVBNkbPbovPE98knPhvmTA5mmd36FPKBg7Ac/ElsvbDZx0hpvfCoK7Ih2zOmHu
AbbUtSyFMgwsHpsXuIgik++JvJCVtiSIS7OsrHTys0aAIM4wFpcMotEwk8Jumf9yYCTi346Xpgxe
NhL2ak/8ytx1TH3TgL10e7Ez4lAzd5QezmsO3IGiOSNP3g5LX8Qyet8DtSvDU2vJ3o8EJprmEmWE
knhXYUfyQ3g6eiiHR7ysBPJJbpoIuatiBWqWnU4jhtiNciC1gJepWtAQsMcPY8/gVJ8DmoHF/yOO
BmlmEIqePedMfBemLsFu7aPEtaZ3XcgIKlZ1aBn+mTPczimE3PLWDxYz77f5WK1BJfAdCrbFPAFQ
yR6nz4YnXcOL9ubq9gQ4hptIv7Uf765MnZB3TIPkL6u++uPSdcXoL+GGm9rN319UCnysI5mY0N8G
uhuDzSWawQPONcRJRrd6gOsDt1z0l6eRhw2wjjfxBAxLFpdbs9SRivyeAmkxpPnggy1z4vO02O+P
DmlGADtzpAeggFdbv/rXPh54Fy5P1VL8BQCeikrbDPCuR7om1Y+8urbTzXx8ZRz9AmSdFrAYEPeL
DtoMoVLQVW4xBJ2FjAPmufR3If0DDvS16q1rg+nYVPuXvwSWCf9cLbvAEcEEMqnMIkTxAVt1lumU
Nr+mGRs8/44oWxBSzDFqJ9yoOM2L604ej8vRQatyjUFKzqZiGUzxX5Uk6GA07qZ12ZplssljDP1y
pvdJpt2DKnLwp6OGRFbRpv90d91idPoPBua+pE+ltOy6/G8Vzw1Tki1S3NKd++faI3ZqKuPrSrhY
SKsS5JkYmwxtjEebc3lbF2I155ghQz1zSDJQludENtHllCcy1ytTu72SgHYCKo4FNa5szWChnNU2
Omp8rjY4No4+OXMzWsjkt1AsVDLffPoiCi8EyxNIQPBdoMF6LGOvJNF5+PwvPITMwXSJfjDGi3I7
hq67HF4i9fBfQqEsX878LzMIoJn9pUzP5Ok8unzKMYFp1aU66EfBVWFgMQMUClcKqSm2IPlT5qD6
TKhk9aRTcMJhe6ckKNd5AtDXSRsoiRnKLpNxh01GT5doJOY7gTSnw1eh2s9pGeI9ZKl1iE2WdaVT
dXM4X++F6OeRw7mST/ombIGk1jNbps4PF0yq9dSh4uCA1g9bMR8wAOQEDf3A17yiP6GTvdvc9aMM
M4lPdeQHF+nH+5fQjo29A6xCRxo3wGSjJAR9v05HBXnN2ukUDWtOeK8h+9qMAMc9LezL1uYhSOHL
zhyGBlitOw0BaueVopCvtEkG4myeYpuRzVlWAXDcdhf1nQJIceGvuRm9ovLaNISXqEdLCKAp3scO
vPNDBNMakUX3PN8AO7evBlm4aRv5TqjuZfuz9aHtw77xIZLuDeJu7CH99CulGjDVXuPLyI9wcopg
Qz3K4pk+w9uNK+hePNCMLLg0Rxd/8cyKl3UI3ufTdc3b4mWzka9ZJxZzYfuwPlKs3Vfz43vNqsg4
6AqLL+vdamc8ItzVANKlMy2kcRuyg+0qa44/wsUcqOUUctPYuUmNhB0V6WuJoQvcacrWl2nGCH7q
JcxApsFfMjo695DMtwkZCUSdarD9blU7hfb0Y5XgOdr6mj09N6VbvNA+LYxFOSEeUhs1+lytLjPH
ODpV2mxfBCUl/WCLWf+byE9iqnGEcsbTdofPQw8p1a38nKB+Axw2q5e+Uo1yzriUpiO1XMiMiy8a
DUchxR9jQLOzkUu68jpg7SnbbDNOGXfNRW4wvfHGMW3L7RJhWsy3UnXfeXI9QbEGZNJu8oaZ7ELU
upl366S1CTte0yZN83z/NwXBmCHie6AuWHBQ07gCa5TFbdPVggqkRn6pMpluzPj9IyNu6gHjYByL
CT2gVoj1ahCnr5k/iAZfszTDLIe5/DNA01oxKnPg5pEaRwiV25sBe2LWyn6s21JsQnwa9hg5S9eX
Nfa6UttS2lbwPysnzH1jqrgy9temruoVVuEygQ90tcJCAVmaQ8fx8R8IWSvqUEYcboCw+3pvgEgt
sMCAfEOMUsw8KZ/3agzr3AATMrXOvMVpppkmEy1hOrTM3R+dmW4C/jV7ZGcPACB6h6/Vv7WvhSjf
AaTOSYmQYAacMrSwqXFCS8nbk8mYQJlS9giKu63cCXB+x6AEEgOmtYrElEfnQE/emhz9OSP8En9a
Y3oGqHsBhCM/T0+GAnxxNjfr0dzP4vue3elU0T7ody4GaKN1wzwfRRkJaejqVlTfHbEUyl/5aAZb
jVAPBiqp0fSQ2JH5Yuwny3JDAmlW+qL0Mtk1sZCIlmh5tKGFFNQ8bmEQ8I5qLJNX/k4FIkUFlKwQ
xyDvK9DHfWrhYSyi/dOD+i1LFlUJrfxtHSCtY2XL5mSgrD1lExEH+3c+vscpTXyhsF8d6fW4qZ2z
728bZvzz1hq1GKf3A04jPefZOZSEAw1WIf26v9gnSNX0eRqbeuuAhXhX7X6+NpKFN8hbFNTiX5Bc
vjzZOeB3Az4qYtZvUa/lSpes82mxjn8Oth2Kb0J9hspsE+up4Yz+7rTSJJA52msZM1MPdOAySa3r
/oZZ4SfOGUkPYca89Eiw0DqxCYDfo2UoG2I0uh2nHQywlyLwHPwcPcKr7Bz3gc0YbFOvV1c0TIYz
/MiTUwHFeiQdz/oe9ArPFoKoBfF2Lsnjbr27QVGsimSvGFOKH6yvD3XCAFF7hm/tWhgEL6JykgTj
PNBfRGLDKKiGjYIhHkzoCadHwUmvLJZ3kOfZYiXPN6fIQxrqmnhM+hbagpyd6SYKEEx2W11cvWxX
F53SjWzIdfbCVxE+5EjfxvCAJqiUV3OKuJAxj+8I2SZAoTOqDQshQcpswkhupQD92uPGJlP10XLL
Kt0x3PAR0EhG1XB+2KjvoTTm7AnGnhdpcPL7g5J3OhdWyK9whC+UfVIhFqbtq5BMFvrQh5dFE1os
vUFJaEfo1HRCuB6psKyE//tzzpTGrnmXKzIFATRgS4YjIvWAdQKFxJ/ejVTRTcN3u8v6C359c+1l
cStr/U+/pAMFO4SnJ+cFGiyXNFmmLgb4msZbXMm9qxpqyh6OelebZBzpu42XpEaSbP52tOqzFy5s
BFIwLLYushb3BgS9IYzX6pYHgG9t5tLrnbYQ7GkkzH+MGfaBw2xHtF0tBdAuFnuvWbWEimm/scVj
/wB6xfX2diDtzbT+/r+LVyDhNhPoh+TGASbIZumb8LxR7eTSTpeJFVwAKpXJtpvaqpvLrEr/HHLy
/QzrgQ3sfyvuFOaiHsly0FZaacITLrgd9D1NYaX3/HYGOFW92LDQZLUjy2DQeducE7sEVRFrzxLU
CyiZQSL2Dq9qkgG/HFDKPp3J5A4wm2LcnIIZgs7DfJZr8cWyyWEob2qzCoK6U7iprei7TsYn95jf
LBK+nRpXjtTihSoOnIPSo0FscToTBlsE6xMrVIw1HS1nwV8T0odqbo0GBdmuroXdtI9zV8o0t2q/
DNo7I+c8p2EVfeenZEIr5dJ9eFjqaQySsHm+t5F/V9EuV7CrsEteyKyPcSlgqLZg5gtlwWgL+Nh0
Tsjuu6yWz50MwLpIeMK6mWRRE0EMbppVTUsjBIl5yLv3Z5RbH3PlvIJDkxtJMRzS4AQ9ecisJAV3
lbXjBAbPlo6BHkXoG7c3cfOYXxCL0hcTsMMYFPoKp/49Wq9YpOpPtznUWef3Xh1MLYbG7LX/I1Pc
5jEfjJvSqhYdntdJJucFJMIU42P64LPlx7jiuYHMwGqajt2xSTv1Es7VVdk05P90wgoxQYJ/gJhZ
XGTg1zEqDBdpfRulKpFfc03FwG6dbsP0b2GIGqSzTExa7BTfUtbjNwtVUtZPZumcVFZPPAe//t8K
LJAfXVpMipmWxKYGw4swQ4TRGu0mbZsBEL8YxZsQWMQVJgRXiFwEA2PxZ5BemreaS34p1YjBs9xw
OH2Bl/M08hIxn83PwHpjrX1SRVHIoyJwm4VoobumhlQyDZx5Pw0DQG/yBo73ZRxv+47ubZwVXM+d
uNh6M6cASiBvhNmuSufJSok/QKdEraalaKD+TaCzZPsUu3bAYJbCAcMBSZ8YCEcsn4EKJZWUuJAK
yS0+OVGGj62kcLHUbowXD3GVoyZlgJUe3lxYY8q1IRjap1GFLdjikKgJsfzbZX4rRkghrUbgE4YD
oDfWnSJVGAIbcs2SBR83gQ+xEyhdO/sIqRFaQyxAErrdWVaAhn/R6SfdkpeC4kx/QWAcviE1BKTz
H6Zg9zQhwJeY0Af6/5Znn2FFR1jw5SnqaYRckmWpdymNrmlAVrP8FBTmZGJXpfwaCIVQMZGpORyl
ICnJMXIzYUd13wHlzFZZhp95eo/6pm/dsX60S+I1zL0ZKOsDJo2n7WnjNDH1ir4kQMbz7sBwhJHj
2HNSnhraocRomNKXnT/UE0ukDevhuFFZRUCQnZqVqVSK2RxMJGuxGCcghFFYJxNt3oB/ehu5ghh4
Qo6s3bv34iNAQjL2yqmx1wpAbNMw7GbL3UGIdPNtaXWdkhDn5tVRP/HAe9OdGDuTYN9i3PYfYWYy
BvtLc3gUwC3R+uFS3EuwQJzl2mWsf1H7yAu0rA7e2dNACHuSmgZ07nyEcNAaP5iemxCR2sJhgQrH
5YFMiJeeWBqpzpc1ILDlKn6siIn3KhV7r+C3uIADHfNipdMspWTXWMqQ+QtcXnwuFHCNQlRqV8dy
xIMUyFFtaEjxzFSFtNhAzirZmWwXb94I1Xrc/ZrScX4ZQ/eFO5aAN01qCNhQAsUXFAA1yCaiLbM3
V9/lZPLh7mwJFSJnXCCI99cQUeccAWlWCX+p+lWE57i9G934Xc4G/c6fM3bRpQ6cEM/zKReptxM6
orQ2Mr689eHL/A9rHmZVj96cXNCvWOKZ36Lk3HBp3KaQHcBLXzzhvK/KaGhEJKy7Xh0EDQhRdkQR
/tnKxP9nn3ERv156ewWrGaWM+Oi1N+UQJxVBLpogvRrcnrkIis3PPepjcXHuJeglhHDne2XieuED
nTEfBJJaMGmqMQ5YkrwJIokLGWOlUrCExJasHYKzLMOdCMYj5OOeoyOSpY1ukMizXVTHKnSHopeL
Z9V53YT2jJt6kfDcWdN/M82TexGGVD81ymSUDNS0pn75qYhcEFPrDsXkP1z8extrveSkRmEwFyXd
yW4iLR0cts6O4TbCjanApxfrMpGVp+aO+qtQU2OdJB265lOAvhO1f/d2zb+M0/XrYFVptXNpKsh1
vs12wCTnc3r6/XjkI4UO+Tsc27fp0TMhrpVYlWNI3CVkmhXsAd/zt92n1h3hI5PUx0W4sQ2vFttK
T0U8L8zGKsfLa8ZSEDgPtmsklg1JdlzxchrLZw7HZlmIHVrAWsoA5dSy87XRET8GZu3PkYyLrPNc
i5Lbm+G5NGQWC+eT5JxP9Xrz6nwGOShgQXhruYuk49IXCyLqA1Cp9mwfg6tH2GNm5yEDQ9NsCSnb
1s5UeXZLwVRSOMYYdvclIrMYciX1Voic4eda7bG8ON3SPnjttyqJe0l9tI5JAjrR4goq8AzoEWID
Chmhtasgtphxv2wgBPIKyc4e7cSS81B/ZHSGA7iqBqDouRxfK9k5thVdAXAIInQOI2X4Rvm8f2vg
ZWhc/r9s779yrcZwunNpzeSVzE1QGAadfhAe8OfSh4fXRCCQNtkx2UzBSo6ABWEpNrHxM9KGI7AF
o2uD6jMqpkjpjrGVaPh+ktf3KEo18ZFXBG4ouq37It/u/Kwtp++8+UbR+/4+t9zsLLGSExoXAf09
xixhDnSm/LmsORgnbz1Ts8zwfxwL8hQReCsHKnFPxhemlm5XVxgO/kIlYFUOkDzNGezONyI2AH5G
bIIjn7NFnaaH/NexYtleaq7IMBpIWZR2bBJ9kM13dHbKzBVh1jLLslvIJfj7pRn/maj71jX3UWaV
ItZJ4t+QVw2VfoLFqCB17Lve6Ivk5LYYh+geNXqndBzuygshv9kOQHryGbD9PxH1YhmQdwWmEWzW
ohm+Mn+SkmNLX18HvrrWOBojfMhFSfPFb3Hm5TMvcl2uFuL/ZfzrTyeb3vq6/4opzdMtnIx5e+gm
ON+UWs4lrG3l0FHEUfV7qYtL8W6pXKZ37WKhCGhFvHlDmPcqi91/jMzZMoCBgzwKDBMvuEWAJiGw
BPCXRAPWNTauUtNQ+wpEQcqJXDG/sZxREynnvCc5vAx6z6IXj2TrqMEnHOODVme8iENQNylRJg1S
k2FB08DhuGU1bPIuy2L9mfrLfCB/qnoRpVt/3k1I1azBP7mamf1l05ftaZTLHsshPGPwk6LsVr0T
lZICPGFitD3YjHHBH9J1RKjPmAxdhBvc2p+Q6ThDKZrfHwJYi1ckvusJX2HUMKqk4Dlnr8dSutqi
1jav5i414aCg7b79cudgROCkBD+3Dv7/oMmOeJVcnkR51hMvfSb3kf34gS0TF81DLMG4BdXDuSGc
76DrMukSuqjpqmMDjspcpjIYqQeQAFIcrvVjxVc+IGdWuPtdeFaLoPSrw2Hj5vKYx+/A+FV5gRzI
9QcbATYIi2G5LOpEz6AnmWPo2K4wSavc0uLW7wh8ynpxRLNh+E/tBSPP+Dzbf6g34Kwf10htND69
VAD+S0caIvTqtEywms0phxlAB0GOR3WY4BBqdUX/vXWeKJ8lSWpg3ImPogWhSuZaezJMwoP8bRHg
QZCs8aWCK9a77Rr6WSne58EF7Xt5gIHr6wZZ30XP7LAu4lA5SL54oPe/UUHRhEbNOOCI+HpTGIKa
+jQhu1PaTkRCydFf7xWs07t9huahNRNp5QvdwgLSht3ArKBViBnMywUYqpWXk6MSe22jQTOtpBoz
DTwHoknEM7lTBCSwpHKeMIhHAOxSYx5qBJDOTK+RVrtZxJwd2Yp3aojmRDJUu7FhkxkMtTWLL783
NpO8QF59IrWqdKN5x7BbPxhwVDNeRysUxahXYkdm4JWiDH/ce5oYATX8muKGqvvj5RLqlApVgL8t
Gdh04GFTveHr1rEpWPKsLtDMhK+qGVre7p6HnxxHl8z82jsQEZ07Ex/3fiTnT9f46GLpv4vjCCKz
qszvDSYzyStYBmnJE0dyMdDhvxc5OM6Q1JkjQ+UQwlfeg0wU/vNRkRFyFY6PESdovUhb8GDk59vF
jC5xPVYv+kWZhW6pk3nyCmgjgfm8wCgCdYI5i8W3JDyQyPMfdHTVZVumIwPnyK7UutSCpLYYRFPB
mNRF8jA6w4p9AIhWdk6mP/afND668uDXpGNTJMIA9SDUNIz6s+GTs18Vnw1uRF9ouwpr7ZTDZxmM
Ukcsbk+bFxn7Ncl4hAMC/wZC+oDDaUrXRBdDoH0/bdFkhExF4Bwc/ylYHLyUSoPcMriIvrU0G+Re
pDK3zWapVCDwOAuETrhZ9TUwr5d5GRiAUfSqu+Ej3etdOd0dAFlbW+ufig00hVZk5ZfwnwJLUt54
+C6FhO7YEuDcQm9OGuWLEhZqepSus4lZLFw5BFcbZqT+GQtz1ZKq+5mHxN8XuOgy5aljV4nHZyKa
bvcqmGqW0S0iEa5e1qf4OBgwjI5Zg4yQ2egXPNLD3s9S51PAeTiMZwt8yPLi9ez3AJuMKI7ImDTg
TbbC96h5R2jcwP0IrWEA1//YqkofhnHZVmbH4C2evLFJCcAzrqD/6gHOyRv+3ilQynMKgTA9t0xU
bn5FXSgq4uMLxatcVJ0wZvZy4b+VAkj+CzXwAOzy7WsMmXbc+XFo7SUREzMeGOEcP9BLeW5rCnvP
Rns8i4VGL03U6vbW++2jPw3n8nRATBLylEtqVaB9BuodgKsnVz+jGysQvJTHyX5mFBPLGVnX1Vi7
gBNbW6DlKBf/RA0czCvulup41T5Yzb8vm1YwohjCFV+uqg5ut6r7bBh52gEvhxbClfE24uvHwuxf
OJh+IKOBThse1pycuoUC3CtppCQ8mje62QtAYBGvHiSNTwfk5ZK6eenM8sUPVj2Y6aRRq8IjlWix
gytgAf6qbLsi6DBnWBL3KZRIsIlXCUPpg9xxpymU7ayJyaB2ABwCmFC1DMCuNHCQaU9GvOYERiD1
ji+X5/mcWNYx9uMBQ9QTq8u7ol+/64/+nRQpaHCqBWloQ4S2GpDwuUhJJiV+sF5LxMlQMm+3cy4V
R8GEN4YPjPYUtNNpQsSffQonNPVAYFOE/4//yoX+3ULBSeOKMZRHeBjy6BM/uKNTmlr6/5lc+t/X
Wv32wiZw30hPLBXI6GHRWbVmtDVl2PRUJCUsoeRrxAWFSY/DC1uUnAs12UNbvdvl+G7DIvnXrGAo
gwQ1tw/pq18dDlIkLsb/9Op6zM1pz+Yh3nS+oUysmgo1lwSef8OmGtrJFRsW8Tbx1glTpZyimfAC
xxE2jY9tooepXA/LPqBicPSbTVEhnyR4NDaaUg3M83WxCmlYlBGoYKE9ZqlFioxbSUCOlr60c/Wk
REk3iWo7JVsknJpbunOp+BSVjpw2KkQ33ELZnoS0gkXohNqMOaqo0+s2I38PsUWdRBI67as/Okfn
eGZXO0zJVRobWtHd21Gr+uqOokEob50Tu8vXBbIgNzItXIdb78EoOq39++yIthOqkH/2+lqzEPdj
IQJIw6z1rytJhScJZQ77Xw7dSzkUS6cl0iPdzjw/dghFAgEJmH6aweF0kzSrb2BPL2ePHtY6p5A+
ys2PTi1KK2tP1pCBB/U636eJaT37cdxdanVPEllkzIesqXE94O3F9y6VWysl6xJ9Mz+Hw/2hp0pI
blSLADAe2gtT4hJ1QiAevCPM77nwH2WvTx9vq47PH2JFX6ksZoSO24Izd55IKQRBSGph1LiZHhNt
4AklvMtG/CyW6+xKRv3WE8Z/qczIXVMZKo32r/mWy9qMj70mkb3/tTCGsmPoB4I/yr4+3CJmOJaO
8ko2z09YToQVxiBUczkJlfp9e1WdhQe8LPOFPuNXrCzauOjcAmBTqkQkXK2hsDLP9ebU2yKnuEv1
9DF9KR7ihE93YN6Ak94ZhoMMLWDAO/y6m0o5G7NXtAKkj8YvB+AUfvm9kSsTcLW7W2R/3Yz34veM
m610jKR0LgmlDY/7ktcjSjuJ/SMhQ0zLlBzNpZDd9MOm/X9kzQq7FE6R/FC7AYdwER8Sk0imJU8G
kzpukFE+DSerahDWd8JP4XWULGmppvWXLl92AIEUZh+Y8+QUCn6RxMw9Vp7q5uppG+UP3fFoBLKb
1zMOppEA9cwDizeEKL0PVII+EVgnDE7ep/6yuSTHmWab0hQtFI5odcPan0MLSZXBDrk8cZH54gmm
1kEJnqkOnLBAgJqOpEM1dXn8F6yYCaKt/kzG4fQidUYqxwwdDjXCp9qoe6Eig5CvZxm2J+lDOzBF
4FgetsgwHdgQkxcWCw0QOofBWo750aoQZqWh2RgPGC4pG0wUIO7fi1eC6oIrd51woCXAVUaCgRkF
NlZqQovM4Zo2MlYsgIZTRlpDs8NFUhEU4cdbAR1I3BjUUhC/OZO6yeuMX7Hymps4TeLQme6J7Iiu
7y5VMV3t8lpRH9MXvekm2p1/25514qMaC9vJ1vMOTpKVYFqHk75xpHHej08LPBSaoyGDCuC8fg6N
IQo+BKhg/PK4/EFbbQMYvt9kyXWR3JYs7/AiD/dAkwkYe7k11fQDYtuVQmksZuvu3J/J9gVKzyPA
2E4qtztWx14UVdAXqNiKzwgN0BDGJV6pAPQScNHpNG+gYDH1KiOUohQ5sVC3x7ckbULjd/jmYwjC
6qyRYkVTXuh927JGFam4V1e8HnlLWFDFmkXWMhpT/bzJihIBvT49SejF7WOhnel/JhsVHANQ9VxP
1ctXnh+QhxDHCxGFoZ/q+ry31OpjDrVDQNyKRRTjO+Z/RDS0kvLLrKt1OuyWJ/zwGEy9CEGc38ce
RvP33pxcT/hdGRFZC2Qdjoo3eE8tJ6Cf5ZcnxEwmtjFy+rO+wIBWRbOeVerMHB/PtGrF1uBTh5Xz
oMhTLnaG8G4RBfMgVOd3a/56cZM5u7+wCX7SATCvydSpdzbxobDrbS25H5NZfzACdP+p3WfszJIU
0rdQkLvCwDXhgiSqXM7XFO1/vfEM0NMPZqg5jrWNadvzBT7d0FpBubheuztAhvgbAMb+zPGn+LiY
s500hBbmUOLRhdbUtvsy7AA1NqzNPOUzVLn1vbcyxDv70F8EjefBSKSjZ/bWLX9hj82hBwwXMEd/
vR7PHMiuMrRXEsdhsnRxu8TjpZ2c2ZdfFa/jmK5mPqzu3BYqcYmkOblDn2KZGe2gab4P4BtjtV+Y
wY2W9Zt3dC7zCmeA6rPySmgJRzt5GuEg9VcTF5UoCBR/zN5hrsb/mLHqGiU/6e7km6+rWdJJ2pXM
RXFtUAwcPsKkURN8mQYLVjbJV2KysFrhJFtn8c8wXW34EFHwgjUhbhcKnKDrU9aNzzpbeKu4hNWQ
BIctMcWnvmGBCsujDcKGRZhw3nL0MJXIpTGd9SyLe0LcCJUL3XWrsv5jZykkLD8G3rfgXubFqItU
aLrZe+HqP5bzi9i4A6uC0Bj7XtMQYksSI0deUTrj52JHbft0kO8XTMs+KSsOz970+Dj9AP/+WHoP
ft7hayulWWb638LVq/HC1XIoIL5JmyUW8ySwIREYmw/HRqanEWSfSXoycaVecm0aFa7XWNS+njPb
7R+fFsoSGckmfnE+YVqJuRlZ/B3qn3SUNeoNgSl7H+NfeCjW+Kgzf0yl9Ax7UmB2/LHNHZCWTZwH
XIIjrPsOgLkJNSU7I4l4WmbEl+Tr8Jqz4WXGhR7MpauDWxDho+F/u01ujv0mmUzXwQXVfRMxjNd2
vKKF39iUp599RyVmBPHTO+YnUere/Plb9qf6k7sFHK8nCpjNpqEyS0H/gckkagfmSjPi9kG9RwP5
WaaqMr9tKOofCRWTdIfOYYC1K3YrvvvscX6n5PWAWKDPT5YYgNYacQYIFLdOvLy2YsuUNnLIDI7V
2Pmev28w8UICN9gQ3m0HssO2lPWrFSH1/jJBAKmvA9pyrbIeeVF/6Czv4C8nImNs4FpCrz6Zveyb
tRAKoSbSDkdBhQjZuXhAm6oFVJKLuNoZV7gteXV+M/DENK8z8vFg+tF97X1QbFOeXjgRsUfOzDlQ
QAxdB7+sCJyC1oEOKgNY9TAqAUllZIqvVu5Gy2h3Mg3TKOw/fLj6qIa9cn2XZRGr0ZmzeH9BuVbx
W9Kg4jhQiCQxUKNO0e6cBponmeErD58gU7PQ68Xyu7Sqfu7ou6HAtjfWSaSgsHeMUe5A0JFiM9vs
8SaqnVlAYBS94VYFlONFWQyP4kXvNy4aVT85crY2cPXQRSk5/RnY2a8QsPj6V6ROPgsdPxRjsZo9
UaSkfJiRSpO5lLQisULfMzIf+kNjjYD7bVnS8HLPEtI6UcYLivS4+SopRlSJiryF7h+zPF4DucF2
3a0oUayjX7Qgf6ppvB+UxXtXdRWL7Dqv/c0b1YbwaCGcc75rRGr8hPIomlQTYCPgL2hk4W+kR5aW
c3erlRgnI4M+Kn50vunrGn+3gukI7l9lNLcWpak8XEjfEwbvUq4/cw/3+tfRP0QnlBElzxOh6Duc
mk7WCSzprSxdUqIwfc2muL0f2PBdBo88BquICukHtt52B8JomCVSlkvrOPVT2j2KBjUrtT+tE/3m
AvcDFeudXDDUwmo+S07R+WUIfn5iH08oxgUb9WDhTP8c+WJnXjC2ZC/ueq1rcf4JVgrwDRy9sLjG
1OQyzJ8fxAMx2yYG3sDyXdEZBJVTq++nU248owx8j0aUDuhoUgz9ky2pa9J9Lb84jFQZY3THLKWC
U6/4yOAcackVYX2kRmrcaO8DNoroNiiZtorDg0t937Jm2itvq1JauOob1qG1YLZiKxUjmNKxsrVh
/+RePr9h2oX1TbqryYP+Nqg7hL1+IT1BVBwuoij1O1D4UCyUBt0VpsEMxtdIGT0NhrzABWWstqS+
unIowAA8FkleSvBD+HBVl3YCYR+wYhsImZ6lo39tRVk7CHFzCNImyudSlqjsyQt8iJYSKY75j4Kt
JZQHo9gjzuO1Xnt+qMRjTALD6sQ3BHaB+NRsTjgWscfaNr1U5o9rbvYhOtAFvIllcDsNUCC3Nhcw
uIJizgJlqaeS559kefScdO7Wfq5w080U8cIkYN3kHPDu8+SmX5B/cuYmcjeCHkGbLZHs3hlQ0HuS
23+d3Zsf1FHjyHwgvS+xGMZYzWQegg187l1w1FZwFNbi0JQOXvtkoO8sIrru+bosrNcnJUck/fGb
GN6aA6Jlsjh/JJ4jcBDDiKgV3D/jbtiojATK7sdUhONqLFXq56V9vdh/4ld2z1cw0Q9zUqsGeoBY
02ba3cMsY0g4q3SdOv6ribDFcBcl+nCxMcKfPuHYh2mtEXS1Y7ZkfjnEFYJndQOM6+dc/A40edrX
UVZVnNwisqcqCpq88q8L54ejCdt8875uYHwUr0cZEaHTVAy1Ik9ubuPZtgC6ViC1j7tm71r0lvqL
++8Wr4DPGecV67irNZSoeWZNY9pKNHDW/8E3uw1LSsfEOZ9H+e7bxMX7X9+r5sKXha5KlMnGMUFI
hBSmMJuO8B0mECEozTP4z8ee3K3u7QpkVAohCaMy4RwryH8A1IIgO6LfNIUHSqueJMCZfCdMbHw2
Hbplb2msd3jkvmleNxzQEXmp8Viqs8sU/vnIoaSMPwtQ7dgCCk4b0AhCt0DQ6SFh4h47AdAsu/zL
xnwOoikY8kbmfkrJMW72wHKp6lblnT8KOBgTW1GCyWd7s9QUGzhJ9QjG0OLJuAxCpUAyLVvAQvAs
xEx576Z8DP5SHBWzvCGquHedaAMSk9iRuY0lDeIqigJQqpnJhwju5dvQHlSwg4d+oCmp1PNY04hI
oHqQVbrwXgaP1u5XlpD8OaBeAvWw9XQlTI92q86qzrzUvtoTL+IL2cdI6uNsMTmVDE+YMDAtr84a
poZ3425Y7fjrp8Q+nIq+ErZuDH6yDYz2I+eOhbkPHBvUk4b1nWj70JRQjUKu/qwzUt7i0UdfQ4Nz
XKX0Gq3hjmLbkbpGk+QmMEHZvZDOCZKGFBflRK7o7nGcq7DWoHaH5ycpFoiitBsKXdpokx34TFX3
WdK3i7HQnQUIyo4R3he9qckQcoQqYdxtBXMaDq3HUoRH0PlZfw+yhrKX9S+kyV9csGGmbq39ehL5
KPwa8FquxgHeBTzdzWLZE9U2OAkCeq+7PiUrXRcLCx/j/zz34FIqBNvURm7u5kiefR6eozFyi0LY
y99IRTBRIqhmX/W04JFdHbPi62w10bBZcmuvR3mikRd51Y/dbnqV+CXJHusBSV5mXhvO8x61n6jW
Kj7WTQoNcoAkhJ+TwPHLv/kbvAlOTonfNUUMApGD0NBrMUJFSWqv+FLq7uczp2ZJ1uYa8sGQpP/J
eiJzETTgq42G41Ff71/XE0P1z0DI7ULwYd4SEW/JzdmYtcBDjBH7Cobp/IajdB/jv7JPwUZTQsPM
Q78dueFc2tGJ8qRwgEWmTnRqUlhl6p5kjIypRHSBf8j8Kw2KT9U25dYjFi5/GSW7CL7EDeRwjFu+
FDcTrPkwbhHh4LGDwIN5itUJ2yMXtlHbBA8zQCkZkbVlcK4e7ZchwgjM2idi1HU5q10R/eWTuQ/z
1W1+NGM78VqBOH+BYD2FHTv/IGzj9UVHKsgV0YklPKBXpZq1WD6oBd252BpkPvGpgeLrzmTLsZrN
2oEJ9neiDW5iisWuNy2FgmsBS3NctzbLNQTaYH1hFEtXELSzUlSGzrspxQ53PWQltu50eur/QywS
kzhERmjlTnuKflKB6ptgAs/8JtpZK+5NoRq09+tZ3clAsFARkhuk5wvODJV+Q1UMG0CxGRblFfMt
QNztaoDHRggn52Pel6D9M8sJasELrTrCisyARKBrrCWSURwHMX4bw/lpBGAp17sLKk5gZ7MxyMyy
p/Ajt4eyC0JZ2atxx7F2AglWOR34k4efnX1z89qiAPPrXaxfTUMOepGPYE06yOhSk/ONzwSiRW5o
H6NaR9MMscTS79kNVF/7OVxSfgWQ+C0teHg1dQhUlA9eki1ya0FKTLaN4YLfjcvyxH9sXL6qLboD
5/XM5Sc+CarK90J5cpyGwZUnKrt/CHnlW+rK9qogJDfDue1s6luUZ0oVfdtpTai2YkaMPJ5Y+CRD
yCs6BaXgS7oWXEeDdPpIpG1NvrS5RmZE+DqsDN1l+si0UgArZhcpoCglUkojsn1wD2K2bodPVfub
GVX2GiQewcl4aIm70n3oSMEBLsujih522iq/TjPZPuvcmvWsqmq2sV5olaH3Z81zlbb7NG986UwY
qaO0Ia8r+FqwqUIYAVoYAY1+GR75PHMIkCiq+OldNSEmxPEvrQldh4/k8Mi7rEV+4bMUxZ+wiZwd
GbIZ5rjoYvMi4jbxeoigaEPvmlFPiQood8bqGeaONKDCeyT8GZp4yN8CpILsCHFEGLuNqKWZwAZ5
X5ytQ8uTr9ZlxfUpW2WW3AWG3yBYN6DWiopUZpf5ABcmKnv5oaUUH7U8AZVT1/hsQczq2xRgqnST
Jp3ibFi/yuplR9567IvbaXd57JMrso1k4cm4vzumu56DNTKT/VQf3vGmeS7rLoA4Fk+sb0i/diNS
Ju7WnNEOQN2OvH7IN4Hl4FeZDf9PTH6MGaXuOUUF9yxThVZe/5iTaKVMCxuMJ+evpPBE4T9okWRu
CUQHTvfeZ3yam5jhKQ21nxSW6rGTxfjaRGfZ0vC0Ah96vpPKenfJRfyF+DXIqf2L69VFvNuq69QH
iZ0HJHJSQUqL4nROIv+gySV5gfNmOY2jepbIBcIRhWpuHekj11ZVRdK0MHedkiT+qqniOzAh4uwX
BCW2vjS3OmxHAXkwgqocRvfGrymN1XWCXRdC8QbBBAmI0L8duUOYXhw0+I3Q0DnKhVs0yAeYZPcL
Y7Y/cfSzIcf9khHCGBFiFytSiCPOKs/ObRYrUAQDgyxtGK+MUBw+S4Q2E+vXYlGzZ64TIX+hp36h
QwWAsloH/7nzsmeVSmyMnTEipSBt54voWRO+1u+lGJc2Advozo3iRk7vc2GEh//pktWshccJXdrp
64PRwQG19f8CCJR8oPoRrkBf8FA/K7xtL9E6uZu0Ml3x/ryOl5yqNgwSFAQzOh8iDy1OegH2rYVE
8WoJznBPyfWC267JPo/cFLsuzUgG92iNpLC1sL74uQk9cOweeqNgZUqGAv7e4i93NKSD273fYMCN
6GC8455l9cSwe+8f0DWBCYDdPQ7G6vOkd4Y39rc3Pp7hisGzXLLhImR8GJEJzRGaPrzfyKqnS34G
5U9z9pyLCq3Byq8Q4txlefgst+O3Y3/8OiAe3ys2jywkj3ClrZflbK6rfb2rXPIf4EBfumOISRUW
kL3s7wa+Hn6JJv4vDCvpDaEPfEuobvDIRsFEhuikNUr5fIU8BAIQJ/kuvBnblACFDViWbkZN3ycy
LS+6qio+KXppVYGkeQPmPOFiVERjpnILwMtuPd05Z4pcdj/zyOwhK7JWdj4H8Hta4hgJgmGAWXVF
+B6HoDdK5EEDD/UCmhr9TVoz8ChJydXAGJQ3ocT1HTLBOktqznt2kUF40y7B95FnJe7+0gr2p+b8
S2UI1eZdQr6ynnwTAMC/tUODYVB8illQ53ShaKD+lGDvaJjo55XMAB5fpbk9tOuxK0k+itqR4NJA
42y8D8S/ycqB6nm3J77W2O0SvBVPBiFL0RUzvwCufa+siLgA0K1kuDZTSS5kwi8Qhuw/jot4CD3h
oeMtmVqOeuAOu4PORM3MCHzp/VbP2gVbc5sMGS+Oi/041dVjxo/FmB6kF73sNnaJ4xP9ToeeKB93
wYvWWpaOMk676YAe/SHgN5Z9WpibuI7JGxI+1LzjV2EkU26AnLcrsltzMq307gaC8hnAgWn4nZD1
h+9GxZt1x/Ihmw21x3EzQW4WYvZL4N9lDRcBVHfqKPHSH9atY5GEzsfE8eQNRN4rpG8LAJfV8Ht3
hJVH/IyJeSSqCHQTplcM3WcCoK53a2paqD2z2Nwi8mu3nwDcim0B7uMO8/Tbu5813Z1OdmMwosY+
NWr+52AVgDB54k1LqBlc8A15QLTFE2yPnU37AEZ3Eb8rgWVoz6+5O8SBFJPpgRN55OMwm6He5SZR
sPjVWXEyN80kG97whf4BZTdGzywqfYepKtF3BovUBQay5X5Gvqt2pwlpiWZTudv16AxYw8nAdZt9
yWD2lNLYK6pjZa759QwTLLuENJNAanri/DeA86DF1Mx1K+MjIRDCR3ZbihdmO4tf0CfPEdoIjIHw
5+udf2ZTf3q1HjcwQLj87XI+8OJ0og0sjO9zb0u1yxKv2M/tjh3KPB+ig8YL1sKvz1018SJcd2Lp
pO1odZ/ww/BaoiiYfAUbsukbWGz+PC7JEb2dx4vnErXwokSKrxIUYuN0Lmn2oPhRgm17dt9zJ9S9
6Bq+TbMHaIc+KQ6Ff3rMruyLRHH/x+nPn6zMpwQQoGj5w/zw/qz0fgNmxg7tiMCpmWScgs4Y/CXv
f8D2c53bkwoXiVv6xDNwJQvVGMnb3w/bFD9+X5LJV7X+0WRdoRKzmgex6DxWjCw6P4gXD0s5nKV/
BbztBewjzMzHB9S2MN5Ms79QNgx7SOkE7KxXccgt5SXoonXCL+rNApcm+iKnupYgtvbqjGpGWZrx
4vOHDDyIhq5k1v5YrUIJHb59vgHXJAHceD7Ff7qU+QydtQXsuQ+EzjvAzr41EMG/GWSvskFwC5JN
OM8/ycNiiU4oBuhhwgD1mPfT9XKJfYViKEWmSos+qULeFQOsVpcn/10fonQAziO0Cg5qhlODVmor
ejjjvnQhtnpriOQ8kEShHh9BrP7oedp42s69Z4EBVATa/c4eS/2ALqbgTuOwQN2bq2mWKloog1UW
S4k+PZMUL/dgXsQm+nXFQPgUdrdgJZihWTjJld+NyJ9MkqI/MOkn5cT/1fahpZzNRJjxzCTlfHws
cdq3l7PYzLxNNWRv9fGuE0gzitlK4B/4KF7Gm0NV6tuUmkOgjxV6UUHaSRq3LTrxmNxVT2P00Sv2
c+RVEoqNEC3TyZQ1ibOPF3UrTUoa0phJdB+XQY7NLZCyrSkuAJFTG8SMUJfxdp+AIeNTrOct6w+j
QP4VVsHcm4VFqAhLrhpo2V1IjKEbiEJeoKpPljq2vVQtwZH+UjchNWBq4q6auR749tFfk9X7++I/
SnbPD0PHQvfqnIqMAGi3pmtZcvFGWJTVcoScgx18KJm3xa+4q0rfa4u7BIcPelDhmLJrDO0D1agR
vSw/c0eAo4My55GLN/1vs2aQN0aV5lAs4gbPkGUJO/MTHqRTzjomLXa3BtIMFnPPpCqrKD9ysmfY
0DSOvLZfwZPT3tphKRKsGwrvmSVD4MhZ2LH9PgGePrxNgxIDfCGArCIPuWlO+Wmbgrv133iRW1CJ
AghkpordXIHz/pHVGnf85Gir/a1yuNi0nNyzi3VzBGIDEBc4CMflziENPY2LiUw5jwbgy26R12/A
jEjxhVpirR5RIc/9yQpcGluC405GiVVPo3vF8x9uL6u83A5nhEw2fRrRI8pRhwhw0HgLDHUrBVPN
vfpxG0ayG/6bxu+pFV1+qOhH1nW2/L4Z8XYe5d6LpBJgwJHE0BMFsTD7WBP5hNKmP4BZ0lS+htYd
N7/7Ox38HH27ZvUfsK51lCoS8uREeh95oMyDqfMq92/8Z+U2apXAgDviXBzWCB22r7lj/pXSzK6/
uz/Vn+rUTdEfoFN/EvnD7aKEG0qhLxCjdanJaCIW1Hy2/OFUEB3+m4Ix/9ccjIHqrkeGiQPNND8U
lKFn1FQwWA9gH0b5uGKuPP+7Gvq+A3IGNcn6DdUL1123dfMMlWyb8dR80xlRlO8WoD57Df/gxqsI
wwBQKNVQVAAzpmxAaBziqW0m8yA2r/TslnK5Qu4/ylGiREgU7EyePgaWvQ7gjiEtAEbRk4+cNCaS
SA6tBGSsthMqxNLOhERpF0y0yDZlcsq1kVgkNLQOYiIgyMFYHTQo5yauFVal3DEfFWc3yF6kL/07
5BPXj5kQSuTBhE+ToixiW5qiL/eOsWjc191z8+Nm834TvSNbplhOpBM+9osgzZbH9FqjGnIFIavD
6AqNExQDvZydGnZ6yA0VbicxKB5qtLP4U3Gt3b7Jfyztx0aVvGBDrDdtbWIdpXbTI0pxEIXE7fCo
36LRw39cVNryGUsmTljEkmMSox2SpX1Vw3QI9KV1rk3vWpnREezdKPc4nd2kjVg/RxhU0QAnrTK7
7YFYLgWhB6aS8E6JOTbt5NqsT1r/mFF4bxdYWW3ycUEozCBfC1gtmR7h/kTiBtNz8YdsmH4bGWe1
R+SKTgIn/+AzMvc2q7zPGZh85vlVV/9XeiAP6SqbjU73Lqwlm5/7XmALHnS5AfU212xmBrOIXyx3
2jlu8EUfcmT5yuBKjnG95ExLQE9pOOxhBEUkzxpRYv+LxASqaTOzeuIfsqBiKEVl708LBUBLAdFk
8qagu/pHlZnCKalHgy8kshpMlZDCT6DQ3+AH9sS/IrmKH44n8HSFXthcqnX75hm5+tQr+AlcoyRK
bPzYNcxI3w2KPkpMfGMfbQWkEnxM9keR41fhqAoddEroScGs28NxJUpJLgkgfrNFfRa7ke9poSPt
UtUAiiNenOkOTuJuS8rXo1O9Ajd0QOTBa7SmrNVpxYAN82u92tu96vM0rRlzrwDXFx2hquCWK32f
iFW/N8iNTGAkGbvG+d1ilMxuBXmTPLZ2K5wZWlGxburYjc20UqvMqrBG63pJhRwzKRG/FONh7q59
qpqyJpxiZzWmd3OhP/BpH1U00CBt4CL5DbSxyKidknlRLNS4iyhManvwt5iLuWEEl47QhyJX4l3d
UY4c2XH21QcCuMUZQri9YcXjwWWeh/OS9tZb2eqkQfpPZvFmtZ/k4ROHTICsABDovEru0HOqMQ2G
Nt2ICbokVETD+i82wyTiXiWlUJYeTlqsN7EXxETSf90Om9y7C4g8hyUulagOAa5wL20VYRdyGSvm
Gb+0k/FkIFrET7y1MmX2O/GaaMh13HdR8wuxFuip4FV9gprYy+u+6Xb6ppCpDgIMUjh4XuYl3Cnm
BiBgO2OCJa8pcqWgxD69TnOjF2/MVLDkD0MKGWdK1c7dilTNdiw7mtCg3T910bypo0D6j92ng1QB
jOGMYko2EZHFxMxmp22oyTmKjR1OnTFKoshIlMNf95rDmyxhVpehfvJEtJdiRdSzXGDlSDaMJlf8
IrCM3SO07c9T5R0f7TGs3+9wAzsx3jb9y5mnvsjhdEIpH1ti0LBNryOsR8Vs4oW/nE1n2ENSywQn
SW7rtjpEWmoOVxWQ4li7jwl20YZp8ofa+2UAkoZ2gcE+Kv3zDCiJiSgaX8574f9rnnqBgOyRSMwh
DjhZ5ZQ9mnPy3whxzVmbetEabe12ifABm2Gr1xz/DqReZAcoZptiiWs4hIImacYKclMwSk03nZ7h
o4yGIzx04WxrLfrE54TqNlwlKjnWQEhxmCdT5G6aDjaCIAu6X1pHy1FfqB2kAy2WvM4CRJ/TfwgA
i2KqRUNrFCI0MIrzGcWOSpn6FDro4PeCIvyr5NabOi6RwTLYjbe2fUUEX6S+6/stL0904xCgq0Fz
GQiPz7Se1q/j6kAPlGdQeE/+1E3SgbBS9UcVmOPOXWddLxHlz+vUvFF2bU2MKl4qZ2rIt2P8EA68
I6zs1VWSxOuWu11jvd5tLK+jBQgGqtkWr4lYzaRFilGuN6N9tBOltpLGQRHo5fBJDJz48ekUBkJI
CRRmWNGI4V95c5qpsRHVJVgzkkdZ/1z4V4vzGpRXIVGkXy77KRZXXl4mce6J0hoIGHaIQiFEwOqV
PH7ToamUkyDM+QwHlKVhvmRwwRIL92hNoykMhJJSm5fVtDaGznTNoZiZz/nHWYLkTwCasGbrZ0e5
fjw9ge3JUTpi94nKTszg00xDv843bd4TrNFO8wDrPCbj7LNPBkhmuhtl3hJKIomsREbn2KZNUnks
cdbLoGygyv6vKvcVmsS7TsiGEmS7UAe07rCBrGatLujHzoWQP3QYiRjKbx8toLpBL9sDK1Gz9mjR
KMA4MyAhu4UYNrhfEdamJGDZFC0NhKXv67Qaw/bUJI/31e/tBpPs1BfyjC6hGgTSm5YpeFgxJozc
sjvVVP/3GrRaXMcuCfIQMaL8SAtl7Uol39K69RVa1Vz9UMpOnjwRHOBPxBH/NLr6UAx+BPGIIf9L
t/MxF+rhOXRlNWS6C+5KGphP/Xri0TvTGotNSmVVyC8g8Igz/fxh1hMOrwcNqwWYsLsGAb1RxIjT
7c/ZSlF1RgCh+BALsg081OzztwBy1S4evhxrfixJzISC2ImbSxD8YjDezo8NplGlrqYej/vdoUIM
HRc7N9qNxVxuiBejNA3MOZqwqDMnIeJMgIRGyTjkgAsLHoR8pHR40TPfjpF/wDV7WPH1UTVftYno
N1l6CW//BeHDj79SxRV2K2tlWknjHNnxSgWwJSu0YxscL+TnAWXCpfyBnbtNONFtbm/v06omEwhE
dTvolnf06i5LIGSi89FGNbjZbG+ELvLQFcbaD6Vy31TqcgRyjOVAoJmQCGfyXuhT6lxVUEZCbKHL
mI+ycC+j8G8DqSVqZyiAIjzAYbWufnRj+QzJAnjb0Cch9jyjfjFe5DRQItl/iVllyK485br01k/k
RHKdTm4dIb8ZFDGYAc/1hIGYDBlzuL2z/7LpFQ1Daiagt4zxpH91spQKPI8Xk+6rBWkzJVMki5KI
Ei1j7ESeU1b6kCxQR3xt9L/rr9j7JaBjl2rjgqUE0QZLAJ5xCmq5MOe61nHU4ULDgwvbinmbGb/1
/hPXm1slVBnPZmIg5FiL8Z3iDgU5wQSs/3infOAM+bAaWBK0aYB1urBBEWvOczbhPAi4K09akOMF
FQ0KCNucrd0AKU/C0hzOhWNrIbI6HVL4eR/NahpDaYHM5T/e8KjAiHMkViCnwrPNd2LzYe0j/62R
IQeJiPvkQVyOKp5Us4KhPkZ+nS7ETshfmiZDSJRQous+KHpktRqCSxn4nI40MxVatyniFinhZxTv
YwDU1qUyMbYG3L2gYGjjCSfKAxBQGefNpYowbUHKALXndag01MHMLlYGYv1kW5QVV4KUGijjFv4x
IuBmXNmfs8Bt+dofo5fZhc7Lxw8Zy1FxOGoehSIelqmGqYE679bpU0bx1zMe/1nfSWT+rRHoR2+T
GphqhZydDFxtkxWdpoq4HdAQG8Ia81aTnj0lF/kzrOOik/UGhnU2ScfQHpmiGv8bu4tcMMB3JRGY
EjAHR3pCvEDpFcdxlDNM6R7UaQguFCa7Xdn7flrX3xwLrA8YCMCrZEGFNXyJyx6DsXa5nITwSupP
fjHxwd1Q8iKRB6PegqWuNNOHrRrJ021YQhbKLxCV7wzNlvgisL1VHPSXloyp7WZMgnWLALjRfZZ/
WzCYYFAz6VZ8VfNTZLA3KlZaasg5TVcsmK7WEDov/foIl0RyWuovLV2cOMZk6CqI+UaRhCYQD8ZZ
/N29gihooRQ9uGlmxOBC+JAK6fUmvtasnrxYT95jnkq6pbGoEWjqnUw0xwDfsqnc4iBoYTZQLrBk
RVYVbc3D3CGhZq+IZ+wBG9ZWMGwhubEL4+DBFH7HOKog76FdB70jRwc1HC4aqaM/6YN3Iu4cv4oh
qbN5FrFTig6Ck8/d6FE7D/SBZU5GizIDQPDJQxGYadNCUx9tN2PJvUf2sriM4AlhQ4vv1c7AoGK4
xigFMvW7N5acgyMl/j1QqjwAGKhWjufmNE2EJ2+4DXjFW9OTCeJ550+t2RhecL2dagpA4XI3LPT3
ocS+rdZpkW9ckgzecztcsqnEjU9dLap+VbZ3ZpVmRXRFN4pTLWwAbh4wQsd0QAoVhjyiPJ8t+RrH
qkUxsczx/LhAouhOK8XgBPqZfaYIdI25e9qElxxjcj4GK+gK0X9OWywvoP05xzAE7cWODYj9NuMv
vsYkxr1l5BM5uwWF7MB0f5lg/HFy/L2tqvwN9tM6AZIVtWHJMbazYmMZlVUPvgdG+iiAsC5+ygQI
w/L5uIW4drOyBRHdykIn+hEX/bA1VuydvqqOOZ1Hi/9TbZCgBE6C+ZOGDi/mtmLW3MNG6eTg8LYk
yAEpSVQAJJZ0hCUu2LS4XuTtqB+V1h1guQKDdQVcqVXv8fr1gPl+BEeTqnSlzJuVmNRoIC9VXT9T
k++LjDDJHnn/1ODMaWlGivMVDmb9lEG+fxD1sh0+IQVPgW0dJDtNbVP9x/uzxD1NDulcfpMAVtR6
QcWtCIOZcXnKY5RWq4TAQSe6R4gQIssFyteY0KYAHauSEveBfhULCoxnwG8kw3Q7d/EsNfPjN8Yo
UOaZNypzeiTkqwocKoJzoD2WGljB71l4JfwnfMMVMrfaRUd5EfHRF38G7pnsev7pArJjzEVbEKlP
73hbaySq1LU+FNPpcfxOQmegUjWap3dxv4ItDkiYwZRlOmXxsebiCK9ismnYVRJkp1YGODJHtzP4
Yefffxyw7mraWcj4mvSHBWS4rqdoZzbhH44XZuuEFM4w7yeRo8PAOz76qYy4GnSwxd6fAkrlbRNE
XNTfgDhAiPcUfEHGmIHdyieq5f5BfVvx5jqmqmJGPRthPJ+SRYC3nTkb7/xTD90Uhv7g1om8+iye
z2vDEVoamhmApU7EAC0+9w1EiaQRbK987RP7Y91ptnKQkHnEd7Ec2Supe3aQDPbjC1lGS1uvp3eN
4cos6C3xmmnftKqD/pNhCeIbfwMaSxC0Yh9LdWYENMdxESUIB0zimGYU3HuG+KSfZ+W1/nBLDTp/
nq6bgvpRRNOHwe4Kj6kwDrS+sWhjXp7sEMBEZoySKGKebsLD2irYUv46Fl/+SyVOG5AWEdS3Y1jS
XjmP9wGVQB/TIu9MhHDFl3J5lN8/jLxKTjZ1qebf75mOWZXA4EeWltjjIj9uu/J2opsdZsDlAQsR
BlXoQSnIcmS6tJyVoDqckBX2yo8X32gx/vTNyD4rFnMAlnmVcljL22fqd38P/dP73+Qr5X8QeMgX
y2d00gtpca965G/xiIgj/U45Bxp3yNfZvv2rsdMvI+aIug+UD6n+d5FXyF+sZZpPWYbjRP3S71ZE
xpR+5sNbBXytvbV0M3xnVD58HDy4FG28465dZNB9/ciSO1kXZ6ekpdvgwB/HCAcV+fbVn0n0Nb5c
UUjXVgxDjUSObc4xU0Avy9Zvk59z2b1mm3BGhiTW6XwuWYFYl4awN713UtgttVirwT3+HT/qsg+M
a3RTxEwIy9pSKy6qJE5HvOPMqJ8gaUWuu8KTnE4sgu+Gu60rmnFK45bBP1dpE8zN4/WT2EVQFjgL
gfhM47d1yngJZnLFT/3vcqPH+oIcdLLKE0MzGbhzc2OkiXmZd1SVYK6V1HzVaXoQ5h3AEoAwOKHl
UQR4iYtCJilKFhwGs2BRqx563MWf2BdYNEEbJEUyu+Ohg7F9cOWhu9dIKP4VDjudbcC1FcImhuJa
76h/LzoecijQbcK0hBIaY7aRYiHMqTU+++YhjDEZ4JQnC+BrD+B5w2uetjYmQj+G5oqAOvDIKqb4
pRziBH7zN0+MXEmgaaloweVRkcVuyysOLZJsnnvq2r2gXsgxZNaCVose7E65+yGR8sLKoXEMbMA5
xij5YqpjuYnqNZskXMTSrg8Dw/X7vcyF/589bYgYwq00U+egPbIqZ3pm47zqVDdlQZgsz8L5iy+X
2hrguPq4hGIUqd307i3gLtW9f0sNnn4dwUnA5he4YB+5mj06I4J0ErWWaGeN2vfSBESnyp5nhAVF
h17RYBqkZf1ZTEIq90EjgJ3u7rWwAs5qJ5r+6Xz1Yp/W6aD2PDv51chQOFORkk0B3Us88iXFfS95
aGBCd/h3wN1GsuIocs87CcbUPGgyCEun2pePOqNQ8Xhyd9IHB7qs+UOFm+YqpQO1NdrBr49OAO4d
JbicQsgStMBkCDpZJoj62KX6N+JaqQt9f/UW5keCC/1PrpCXm5ZvM2z+0hTCnHUO1fUkD9EketoG
6pfAE+cqpVk66ocl8e4A4EKuJvpQ9HiWV+va788PdVKEN/wiXbTf/TJNqKktNI3ES+0eHTt0cPoq
oeRbc7CImybW8GoK6avPOUCfewk62k6jlQx/JH40ORez3f1D7/Beqt1BcaVL5dTwwlQCLUoTrOq9
FXK/CRHACqKL1XGi7AvKfG1mSCwfZ5/jV90x912sxmBSxswaunl5j8EuedtG+npoSEUoCIgbrjs0
ZClyAJQspgow6Id0J4q375DD/Cm0oYVauz1wM0UX/DUujXHhIB5wpvcb0F07JSnPHcK69e4zCBfD
nMLzmz7xDamnpowFa1d/v6lxFaxFe/9Wc9o8KEtdqZ9oOeyUnGDio0txhh0lOJZckl0GHRm6Anau
QtuFCopBjLy74hk1y/NTkDHaj5Cr5XEOLwEtavw5iZ+lM3eBWQgVBqK+OhOBflkfWOfrWcksAPtL
ji50ghXaydYSr3ipTrJ7xg6Qd/JL2qMGoBO7gNWXbSfHthXuDNbXRWIt3D0zhAaROnFv3AMTKFhR
AIAYJlB/TCABqbtYzKnzSS30gtiwCcbI4J+sLK0kkjhZN99H1m8Af1YqQ9AIEJoZq3UpN3+RCiAm
RUjFwzD8vI1cyW0doBgzN4oiYbTWX1o723Yi3stz7rXgkLvmozVdcI0WUJRrbuKTu1EKqfT0/sHs
Jl2Q5jy+7vEalC4uXQW7Rb+MsqvBjPh5456oEJOoA1vt8k3b46o3y7eKmTjm8KOEjKWM5PuNzn7K
t8CLihe00nsk3OHpzIkRK4YhQPPd0Z514Arha8rZB++CrIi9CYsg971LOkmXMIMcQNyM/E+y0Ak9
0PNPkBuq1p0cA16lvJDVadUHSEEKl5p8GsR6X+swhbi8kgddX2UUf/p4LO+b14dMcq+ZkWtXpjkZ
gB/TMkguAfRKBEeiiebjAsPdAQHDbXIHC1SyPojIfL1A14Wmg6W4emVyr1R4TQHoIFFrfk4NtlN/
P4rfol4ejhobGiiGxzfUaqJ020C7XH5hDcF9wv802OfYcSnPTKw7AewHP6XVZPlEcD8mjuT46EWr
V7fjeKMUuJj/Xb832l+OjZWm4qtlk8zalgTQeMsJYk3oQz9v726sfOHnCix0ewzj72urq4Dt3LWe
puf+lRNauiJ3Jrljowrok5wM3WJaGrakV3siiL1+3HfR5CSj5iUv2n7UrN0vjBC7oDSbupJ3OFcw
VXtFqAtQucPYyw3h/FVNSWpF2C75dHrdgfwehzVvV/MU6l6va3fJ1SsHCSRjoqWo2YUGYsEYDz+z
roCEODdbcxfIsSsTQSAhLuxzw3ZXC+VYWlgBowdAGBjrDMT3x5NcWtARxrxzxeChFXDgm/e3mGVm
JPpNyOsWhjiophtzAc8FpLHl13g9nGzCEGVGBQWZhLnokY1j/ru/xWd6FVlb7HUhgA40K4dpkLnW
4uGQuDC4VPXqRQ5ACzcFFSJ/zCbUdvnWTT81U+CqMbcpsEnYSWaN4+MYhfG9JXxpZ0IwXp52Kqfg
OJrcTthLjOB0/DVGcUZguRNDfakBNRIFxgQGtDVSI/nu8jATJMh8KVQajh0lIsbiOn06i8gF4TYN
lVMgMv3OYPcjcPlzsaX4dfU+/WEv0H9EVLJOptZxheANB2LpWvojN5yg9sKrSEvrUlMtcwcYX4kQ
TNEDUOcmGo7pJY/UbCasIxXk4853LjZMWEaQD/KWF75rSrI4ERLY8C0q+xBKyEcRaA7o31R2srOk
QrMxhR8h4vtKlp9GYyjZzJhEK7S0DKvxMa1YKXZ6L9+OmqDhC1onlWuH2qLEz7fZISm05zVedEq0
F4AyehQiww1hFPYUw6O+CqdivMx0RDC0xyTJUNLh4bE1ccinq2BRGYx6a4dsd5o9lK7zy11dUikE
p1K3WC2RMMXcRnuRCzBBa2twUvBrOw0h20ALod0KNVJq2PihA83qXHoq6H/l+q4wXL7SnC8FtrVq
/5Ru7CMKLi9UEmlzBUm8mziC3KlEZwrhf+88J3V/phOaShQoJWZB0XvexLTjXuJ1rkQNytAwgOim
cAFLh2VikJ1x2di0lCjKSoMBcQqA8P11uW8AeLykDPNsn22HtfZwMmkuPUUqiID/HyhTsZkMcJNv
W91QFE+UEDFzTZW0cBaKWvIBbqau+W6PdygLVsnhkBDbH0k4M7xVZG1Ph56d0BPoQFKZc1BYPSpM
oqlJh5nXy+Tv/AsmMHTd1YMQhibLrUBk2DMVUK6euUe//h9YxSNB01aKZTFIQWVgXVhcq1XkpElw
PUXxRVSYp3zEio83MpFPQWqu61edYrm38LwcGfTnA1eOt/4iDHgw1Mb54/kmBeH5pBM5RS54IUkh
B1T7B/kQIYlO5e79MhtADrAWqQuxH9UhaJp1HiYJiBkwDmytbYmeFo44LUS4CUrH9PZezarAmxqS
4hro5ACdbt8ISOjmBdGzeNE8Ve/tc+BSZbid2L/rac5jLRYzZu8pMXBW/QsM7BfdZ/XDOEQ29u2Y
0zd1MVzE/C/6RWge7le5HXbghgYyZ+STR03UiW/9UOTwqGrmM4dh01l5GM/CJWoQKrDaKOqQ/ETO
2T/qTvKE11Svx/lOsQqEp5M06ln7Labs4rfPMONDdPty/wgtm+WZBryrLiysBKM30tbnloMJuJ1s
M5ml1gv+BZfoC+czTyQab+PRJWfh3QWnpV2TJSnmGbt37vTdTpiFFeRQpMGy/Wbae5v9/dh05J/7
x0Tvwx5cfvmX/AIViFdUHa8x+NWEVoZ35185ghiR25FBXpAcW28j9b+k4mevIZy70Jgv0xBpHFMZ
XPBkiz5NtYqDqkxNrCOL3FiNJTs9qblbLqNfFMUBftwg6x+qOWexpvnRodNr8ejEoD9OnRHWdOjk
YE1IaDM2MpjQNABuqK5aoHgv5j4ywiDCh9oNRohAsP9goPVg4QhZsiuL74UJ6NP5KDs1ID5JIty8
R5i4EnYR7ktG807QHaGbxDqeQVtEfksUQJmvmw5+EERTyQwLaOLp8riIjAHhPpZTSuXhLgit1g2X
TxKqFxgVtV+/y7tMsIa+ARKx/7+pzt2RLSLrznDUrltBWZmnAKjU9jBDc1jNoG6OHw+gxIBG3lwZ
mTapDY28v+o8f8gqsEgoEAq1el4FwuP0Cal9XwwykHS7WqIkshX4yAQg6kSObja0O1lBC7euKU3Q
afSkR4/K/aUNEFZZUdJJU7dOaT5/BV5zErDVI+kjeX477sc67iqz++aQYNSyoWjtdLQ5YR9cWI77
/w0zcvAXunEnA+xMgUIVPEqySlTq6vLPgISe283Sd6lFez1ro3GAycgPWl3N3aVgzeQ+uYTo8Dgw
tPiSIrwQyaFOF5hKTlqX7DQynoJzCVN6hHm+AhUgkkSrOO3FCerrKKVys/YnNgsukc6p+Yn4B7jP
cUU+myudcWvvijYiSku8yc5rQarKFktcs2E1FeJNfigPbnAd3txDq4FiksBWppjj+/fEAy42W1i+
325qAt+Oe0rzU2sfJJD8PABGSbBS/1PYYugMmEURmgrXRNwXC10iZDvoY5M61r+BGv8JWx8emG8P
KjTdUGpzBChcchH40bJzQg2nFRgxjtXprOSsdGJNOAO2F5QqZ/UNMwSx0uh5aRqpsGbkIInornXZ
nXQPDS6BCyujqBANRGTALz2Y9w1KuUzCtS+9XZm2iDlHPazxFdV0eBQJcLOhEGbP16Kl5rNWOdXd
IR2q2j4aW8iRhitGLnabtXe8cc6YOjCL0TYj2VXTYGMtrG/uczD/qZFjUqIsVxLAqVJCiKyal9Qh
LSjY5vEpWm67ZCP3t89dKpLmMudclXgEtHyy/lStgw/ljL6Kc153dQ1LiuTdLoXnvEwNoXaypeUn
neS5h1+/rIGa5ArS+GDL+a//zXlYogxf4O/HYk5BvZEeWAZEmKehiZzP+AbTXLehcYZhBx6oP85g
CgrR4PDOP8nnQ5f+nYRFq2SFrcN6z24XRb4htialdwsU1bNCCvgJpo2zx5H+TcpunRqfmfzaJ/jz
5qUx/+XPK/Bq7zvj6nOZecfCZ2+w7V/tBJBiK7Vt23x89ue7eWpNZzptmugXTCcJ+29nTBFF+lB8
Cyg64Zi3bkYrGgQ98aL4aRi5BHq3qIa4LcJYftTmXa26ZdWgzAOxCY4uuu7ENzzLK856UEoY3p75
yIrNHI1Y2EHIAy7gHYezXhBQUULA1rIpwGgGyxetJFZbaheWb2xu6TJnbrWN+xSHUHJ5xtvG750B
fV32ejejUMMquIt6fsce3oEnG6XOpIlD3xEmOQD6CtKWgzwi2+mBgytX44/6bUkPotEKhTVMIfBS
p7jAvu2Luu+Mg3krJNHYS9MaCW8uqDrGQfxB7K36Own/HPZq88+sLvfnZg1Y9s3A3r6TAXA9QUwR
xngYepNQMHpLy1hWMa//IpBQ/wlygu+wyhOqSP5+gH4cDMBKunwNV35A83i1fjJGEKeN1ArYkL2p
dlNyFbPqUbkNVy5sNmAM6om60WswcC1wvDaEF+uQkoLbARk1qq32sXlwDQqA+VPH6Lb/PsepMkom
OvVoOaiq4NSDwqBfxdIj+BzfoN4pS5n+mMiHjOTsED2SkG6CRqz+1CbxJkzGybFpgW9sSGjuF2Vf
X+jJt9Wkbu9N6B8Xly7n6vD96qseAOV5Q0/PjkDTo/EFONidU8wQjti5J5+iRrUfSHZQd0UfS6uQ
NAbf3UVtxGne3iF7v4IuSsqaP9vW3vrID4bzZ6t5oDRxPBjCh83a/6Ot94lzu6Dn7jIGMmc24IZc
YCjyt3P0Il4b9ymQLNWqGNKTIZ3Ege3vOaHHp/bxgcy4abythGgzbSBxhgg+xtFmsloE1kV67M9t
mYFQqyJn6XDxzD9SEIVvUDfJPSwxw+4RDSPxnsTWZLLmRHcBXKrFZTtTuSmw8mOqREDZoFrhc9AB
ta7ANU0/ug4HppVYGqcNVEES36wXFQhatmm/JIOh249Hpg9a9tSpN7RSArE3akSKKBFGeN3+6K9K
CjvRjFMZJ2smWxVBfXrf8J6wvoE9vO+jdwcvtWEw3ICFeUscxsWRnk/6Pzy0O/QhLoHzNgSSZSTx
mez2K473I2YQxgm4wpPHHR0v973tgeh2rE1bBnC8oOaxaxp+J6V6oMjcRrw3/kWC64L8m8Dp/D08
K3mruXUA9cRhmoP+p/PwQa5kBY9/H6oVC+C13LRanXcWX6qJhCfTs83rN8s2iohhxaIrbWzaPIGy
FczyImedDKAJ/AfYBSnuHJc/P4bopmkUz+WDPv9GzkZkMusfnWNVJ3ogNN43gcMeRk/F/8fMzhSC
M4zFxRy9ZPiDlqJtSdkGWVabp1D1wrh0Ny1eBOE+BkIH6HKyi4wHi6J9Q/plY7yJ4PtWBbjSlRRQ
VZaRCGp80iZcw9DaW38Up7d8oHvZiZuUQPnai4opA/LAQPqBjM4jZo1B91CiGkMzAqr6R0UUJ/hG
70zYE2oeQiq5lUe6oWhrKlk20eAeYhjNm2Wr6Z7mZoHJgkcnws0Ib0k3ujvQNycuian6XgH2bYVS
wpwE+hIhQwqsuseLdaHJ/u75A8seZ6jSZRWkmiU/Jd7OjbYSVgsBaxhff1E71hJ30swgTGlc6X9x
3I1ELmxbuKPv58Kw5Bx+iIMm8L9oZB+EA0SZqWkTfZCprh/1Q9rK9u8qBeDtvJxItOe/ldhI02J7
MCuhm4DwmOSx4zDmO56jXlM/qbw7SMhEQupuF31UpSOh0DVTbxDNqjElalf7CNEomsLLXPfXQu95
/iwOXsDoeFnB3uORifALRb+AP9y1xxRzeiZyJ5l1C+K/xOcfzRuDg9hgqHvPUdZ3+tQM+4qivUNy
BaumKLUxVzIUNSXTlkU+xWFIAkZKO3LGlX+5zu6zZV50j6vkAnosbo21g5gMfNcs9m/bKF9/SyZ0
eDCFVWMoThHjE430J2IMfJ9AMxlupM+DttE8VH06yu01epWd+e8beAltFrDTLNyj9GMvV6OZTnTx
1CsMYfuuhnxQBqKvPvoZEoG3TFusg6XQVb+nC0US1YxmlxYGuRX4DnZqEBUPKWdpwPJInAZVnlpR
bDcnwOtVTXGnGWYsMUEmYkYXaFGbY6L5fj39WTlCACBVigvHNPLKsvnHKLGSkJeVLLO59YeEXu3B
pQfDhdqh6iNr5oUEfN/aK0pl1OGtBiClkwkxicRHBmNKZ9BcmOyWF1H394g8mGvN4Qtf3QNPpMtX
r1QBJSFkH9yyxUCTmLQH0wThtbcueegQ9Div6yoM8PnsVfKZc2mlSxAdDeDEavYhDgK336KtpXRR
FKhJpetIW0TXJn6nrGKVV8GdTtytjQVoekK/0B4DhH2ZiMjUz+2MatY6jZpblSDc5WGVWLMOLFn3
CALT18qlfBWv+JUxG7vTgh0lz7FsJYpbuy5nb2wfr0TyDFxkFS2Op85aWw47tTT/0qlWon1ttx0l
6dYlsp5VZD1xakxaUxBALkx0ciXxuchbL4Tv4s/PZ+ubOTo6oFt0wwS/IypmiMtlNyhBqBCzDgsu
qlaMBciITbrA5EsRn2kA7IV2r7BI4/ALS8cil5UDUyHGvqfd4fQG3qz9kywybkkeWXaIJi8P3FZH
5KM0Vl94sDPSgGZaOzymAc/Z8hBOAWazPaosYNZfwVjYwuoUPysA7zZQLn4OjoMjjATPhGbk4gB+
7BkSVfFOgGu2Kbo+yxJyfd+ieyD8LVzLC4+Sdl+FfqRepNAHWMtZCiRHPJuc3vzm/3Po6KV8RO/i
NHyGiwFJMU5MvV0DhiCphtRs4gWBxRvfqm8uP4uu5UxQKqBjO+2xas0Txk1lhcekwDMJPpctWeWv
Ml8GQcIv8vq7qOWEW3pI7jmjymHkGsh1yjDBNNySxVwfCcq708n4R3iqdHXq8QetPb5hnTO6Unpa
vdTfLP+PnkqxuwHrs3AG3SguvFyn6gP+Zp/uvUp6rJkQ2nnfZwi4CNOt/hsK3lnQ7RRoFYoJmKr2
m4NXeB6X7hZ3tAjWYln/SR0TuSZHHzL9JlU0PvNoxfnRVt6uHOigzasPxeRIMMuo6yILldwBWy9W
nx7GBjQqNGxITKm7jH0iUu7p5LYILFJrK4SQGHZIV0vKY1KN21XkWHADyXLyJ3S0cXw0ga6rVRhY
qFXAAurVOkUgXOX/XnCBbkB0rlNVa97v3hv/4ZonNoTTDVEALeKze5JArkVqqn31MdGQW+x34mq0
ysij2jrmi2EGzU4uobQS2F3n8OpOLPw1a7VfaOiL0voI1HGcCDGKYloJYTPA8W6YqfgLfEC8qwab
jltymtkS7mKuqQ2g2LXN+lQ/0rlLHg6magEE/ggo+owL4xnqLvSfUxejszz54sNgxc64J0tTvrZp
3SWTOGXg03Ri7jLLjWeU2aYklJy1KlvpxNBcwTHTxdkXwX+3ME8Ir+a2pigygQsnbwBVXIkjTreV
7pIK8wmrXC8XDEdiQyWzFgVyjEFABC21NQiugZokbnfolLqLBaOCVrBATeRONxH+jhbUpYKX2iBa
b9rfyOjVDGUaSJ8vr0v3QaK6/6bDxAu65tNuFSJpFkfONhrXqR3Zh2uSAEF73OWZtf3WUvcRryS9
WLG0FkxeU2vEf5l5GKwozAud2Bkv9ouHS/CBtZf5ZvqdPBM4F8rdQxyjWGzv4BfRGORLm2qjUEKL
+Lcy75VDpv4YqcJiZuettXKslpEx4v3Muoql6wOuSPW9zOJ3L/vVmhGQ4IkXBNrKy/WJwz7JkOaq
OTrGKJa9AkVBXkeyhDhD8e9wko6c955qLPw8EiELuKD2mBcc9bxqLLncYM/sfVPBk5oSbnj2yRaO
d3GJhY8pS7vsV5NMnSoaHmGaipduV6olQxoqMTUU9aoC+pu8/7wwed2CYI/zgpwXQiSkIqM7SWGS
OiTgpM1Jxn1UkmTrabJoT2b87mt0m3tRls0TedBt0IzYU1ta3PSdg/iZRFoeOQdBjaCE+PdaiM99
DC1ODqVFtLyqiN7al18+Rezq03yBcmSfTJgmA/myi8tioRe5dspNMhLG96dmEb+ZfrvJHIpSu66i
cujjTBlrMBoQ/+wnWaAqQLmrl8ZOTlPGyUZ2Of1bV+FRIIO+7VlRBmuDkg7UZtj9yRpAbUrTvujz
iazLYgG6dECpVEsDnPDpM2JAMgMIySJOZZ+kPqp+EURpb/hPN933GJYv+bIoPOfwDe8fjwIGcSXh
PPMXAjteiuC6NcF3eAbsEj9J+UIKiCD3rvDSxKerRt+8za1bLpDiKJr19eV5HgNMY2u2BHsiAdVS
4thsKziyAHebUb4Skk/A7HGFbn7PW064A3zL0ftXmfrqrvEXvFLuaLvyO0o5uVirDPLx6/QdFz4k
mB1t3MfBg4jq9sBFvhex9RhX+2r0y0sJzc1rmUqHNHYffnYCShGo3kH6xbKGDRedF/xMBpWGWQxW
T4N4x6XEwcEaIKV5dSCIPPAJuHIbXLi5/Ms4Ab+NaHCAX/RevmXsAIXGejZd3ecWP2TLkiUaAYqF
lQRn5SHW0iv0UL7tPY3EtvXc3qisqOkkyVhj6q/Fo18pINCIGfZqxFR+m7k8iiTfPSurQDR9QlfX
XY6kJhGJQCEl72khx7Pkyy3nuQiAx7d8HHax6s/wJd9k2eaTVJz4aIApHoll3FqKXzU1YTfREto/
VU/QJ9K52ebLvHQz1URYX0eLdPQSJubBIOr79x0DFsniWhN3CycG5jf9YiqGun6CsXLTyDm8wD66
2fywaDLbRGgImVebQTrAmbFsL3Yamejimay3LXQniiWxk425miLOD4xAeoKyBQTXrJTZN+CSnZ8a
lVDmWWGZCwdDOoavfvbxQgS+pgLTwgX27fN92OIMz/uDHkkjA3Dj9P/QW3XSd3A05UlCE5H2ps8X
9ufzTMpbG5eTixgAsbMtnwRM0NcMFgS1EKXAmACzcx2NlCkZP8kD/ZtHqB+HdSBMo1suyBm45Dw0
Sv+Hgbkjl3T+vvlde/mPKmjauIrm13p5EV/gDzyStwq0FSwHvfbyHIB/dejXPjD5/Hdx0YPpQjSt
6+M8Rzq0DIQewu+cEVfvfY1u16nsmvQTQ9KvwkDxjPFQKSGSf55XtrXjEw4vU+WMLiCC2eNb/6v2
ViMVZISzC7BJB4SNWtgXSBIxmrgvmZznaUAlcHRuDUJb4vU42lH3fDhvyRYDIFMBkrXq0vLzL1xd
I1NkDHk80bljUf+Mpz9mVcBjbWh5DL8R63ik8cZkbp8GfVWTjQRCqViv8jOfP7zS6pg9COPE2D3m
1gwFN/+o8r49y5uD5EOX/uLkB++v1/f1lFdUAavkTXDHEvqBsfAMy08HEvipn8W+tQX9i466SC/I
jMA087m4Da+rTvxh8wmJcSCWLncC98U/1NocmYcW9txPPDqCeGRcO2SpQG7r20N+u7Fpl+zyMh2x
XVl4krcRcLWHuzdmBqf/rTuwJu8q2zQkMnqBqNtY2m9sfKh9M614/T7ZKU2VUdjLiS7tNcP7wSHG
1LO4nrMGneXQwPiz9P9dG4fittqpflhSvSLcExh921T7Wl11hyk6rk39EEPNY10Bzllb1/IhNCjS
AmSY6bO02hwJhXHTgZZqTdP0N2YfPLc1ATLgk3wkTZSvStQhjbj9AHzUEiUXG4CK4uoPsilpPhtS
uFHkh3vHA5s9fewro57dK6rFGMGQCTGhQLE62gwftc5vOdN4++AJHwX10vMGI3o7F8TcbY3HmbV4
st2ZxzrUYYtZVdVip9nuCK6ojD/7R45IMZQsavmZWUYr1ZWbG5SMjDBjyIqL19fPZu/y9mKwGNew
nzWUq2nn/7sKk4x4RzZAbFn8/jFwa5alq+JxEcdg4GL3wZ7Hfm6Wq96arAFLiWxqYlNOE0dEhvta
dXR47wfcRd8j7tCtuvpPso/VqJUBGR1/KF0s3qtpz0TYT5VVrM+psLp8z5jcmq/LA+6+FUq8LUtI
Ox2c7XyqvfWGCWOK6KCFQTv826lIJjkvtHdf/uOWGwzLYtmQ/KdZjKTLJC1if1dcvJXVeiSs//Fh
9hOwvdw2KWnNXDL5Z9yg7duHEbD5CaoQ6JHRCzJimlUDxn80IszKDGC1Y1+EDKM9SSZwbkOIREGT
qyqefdKqRO9jXQRTE7fH2IwBxirSautugMoIs/Kt3n7QZumIRBKHTKKoJM8TlBCTEU4gMq8og48H
vOE5J6w8DU8jdL2XGBvwn1lDnYxvfcVUuraQd7Jz37FEtSsscYKaGjdXvElEPtQUIi8lW6NWOXHi
Ftu6itGwYsKXHoQ4Yp9WRFMpY7G/zjf28fzhrxGeJAcZ1K30OKgpf9IoUwDdqW5xAvK9/suS5F9c
rIWN2DmX+I6A95QrCk553R2rXdJb/8sUcEdl8gbXf+ff03jjAI/BdDbtilBNbSSm4SK8quzfnWnZ
49qXlpJ2cBx7PKRR7G5x6VNcgSwwkeXrnCu4xchmARM3slISfFWvad7AdQTQXxtDZt7T77zRulDJ
Pdm1LyyTCXk6HwduD0QA/0riuPVsBKEtLFsLk6U1qXG5QPytLp6IihtpfJjxgj636jJ8Mj126Phy
2HTKtVTq+mEKrnBsI9KBGtNygQFCEb4Fk7iSeYGI5+YXDobdQPxsXVUtmcyKf1XPw/jFtslFkTwl
Vma83DHJFCIMvXehJXCQPo+OPf5u2DYR4iZFI2LV7GNAb0gth5+lDyrhknISQtTBZzXzIntb27T7
cCMB7/VVz/VDOzITOInZVppX9Xu1fVvJ72GaP2QZUiji8j9Nd2vImlJErL8sLBLQrZwTW1MexWMx
z5D9TDY3epS+CGZAGwC1+sh5ZJsyPxJm6DzE8jADlRj92qMt2WV85z+QjssQYLpFzmR1EBRflJ6m
8Ow0wwVpxR3olCkWdqEGWWL5PqHvtoSxFUcz9A4SgqTITqgIq2EZLeHFixUJrVuUgfYRtf3ZaX/R
Ebnuvbi9TOVR0AN7yKmTwmXLWR387+kBdgBMluO8PzXNhsUjW243h0lblxp/JNHDcHnCi75u9Ehe
Fej8qKOyLGLsjxZUqk+f+u37r3wTK3OrNZ0rwI8PjI0YvZhzuBPBXqri3R0mX1dCm1CLtaVnkoEh
Dxl+4FTzz+fG5cP/VkNEc2iewQUW+b3/EX3sfvsImI/lKXtTYpF8nokgegd1IGQ8a2gF3TkznePg
xoF0XhZKC9rqPlNORSaG7rM+/0Gej8mTvyMfpdcbZnsAt/vSycWw4PitJPRA83fFuBujUfEtmitQ
WUNbE22+2NEyHXCp3KpR1/PMUUa4mi5fO8Ktyz3iQct4b96u9siF/6s2G0X1AeTFaeqzzMulIhKG
ci2UX0UMVuuK2Y3Z2qI8YTA2qkqIMU5K0QUthUlqptmm4AQgctl5NAfCbFmToaWirPlXwamu6Goc
6T9FwGLuZPYTmwWo1zPBWnABcW2GvAEW3OQzfBQamppK755pYeTso+O54s+0b9SwKgZ0SG7GrKNs
mMy9UV5+Jo8F6RVGKBlgq4621i+xDfxscgxvU6iMHrE1aEAHe+Mmbl1SowhWp0FgFIN71Vnn57D7
puwHMQ5HQKG6yUw9AP9s6TWI6FO5mgVMPE51q4Az1nn9oe2SD1wMwQVa8TXHeOux/ZBYAAzH7lLl
9xBYm5U35049T1f1o4UADKcx4ORWmqrnMn59NE7THdKJ5sWfT9tkSDxhG2p8mz3Y0XR0lwbLYvBC
nJOfjiQzM2QDuugZ9jAnNaCD9jfyw7yf//vliJXB8bv19Sb9O2gd5h37IB2Aznxr0it2Y4yXMObi
WRMxUQYrg7wpRcurpGebNVIwxagmAEKYEOzZXXmyi3aja4FtIdiycrwlWKqCY+iMaOh2F+gFyzrN
0sXC+EV9V0Kw8q2QAWki669oGyDGlCicvpc2fkjKaBQ6oQF2klUoNoGThf0msnGj+qtyedFnhuVt
IOHekuM+07qDetjsOLCLkoKMmeoD0IxCDkW4X5l7bsY3cHyK2kE6k9vOCx77zhvetqoMNwBgm2CB
LVsJxmyKICObXhM+UoYj/U2bPUwaORbuNg61kvNFkLRYfp0+n/9Niu7zdgKJyNCNrD73YL8QRfft
clz3IyRk+wqI2yBRclhBYRjBKofAsdpxSrKhg4q230L2C4eAa0ny4r0KKeil0Au0BHglOdFmPvzz
xtV3c5R7eDt07mA0Do8jQZe1mtkYxln6faDzMKg+MPoxKCjHeeIB/JG2xV/raV+r7XFYNTBMihtb
+ECXo3whcXjjmZxwhxwR50R9En0FPSuh5oyQorBU8MKMRQC2rn5PZnrYwTbD0gJT3P6G/IDsV2lF
jMLC4KtL6Ixbu5HUOBodyPn6uYPknxVY8fP07pxcq4JlYCBQpEjC3N5QaAtI+JPxKqAyM7d96qHk
G/3tGHepSoPQH4c/KIUj9E7W6clRTK6Hb0Khk8Ty6QCq/++ngUq1ZDpHlEoMAdQE1mqQFqRNNw0z
HwHXRTgVd7NNXBreb0ecfMB62RRbbVp+Txl7sQJJhpIanj4YRFEHsBCmMucuaKPVoVmPLkNL0TBR
/gKYptSF77qmoNTjAP40Nz+WoZQjLgVlT0yMs2PkCPFjnWfLBjT2OJovXw21pWFdq60Zsf6TSb5d
FhLy16S35mF9KYEnMQ7IGdbqGv3dLK8VjQpWMo9HEP8xtyEDhdXA3GQ0+9+00zfJpePUhq+tiIeA
dqEsDDJBrelc015dW1gh3HhStON61WKTu1GBKdE64ivijT23T852smQcQzCroq7EoCVT1sX6yTQg
YaZugoGY0ucybL9CXZqUd5dpf7KEcjroQ8GV5WXNalGhwJYafMkjPf73JuJxBX36axaJraqAjd6J
cV53KuTi5VB5pcSZICWjdR2e7xapwYH/hC4zM14Zmlko4dlC8QIpd2K35xWBWzMdJW4c6IkW3Qkp
WN4HqresobFEn823ygiimZZv3i3gngpU8tQbpCdFnUKyLSDovL7hljs+HslZwnBMut5Nj2kE0AOJ
7ydfg+ZU6Lldjl0LX4r+eI/C0owKV69gIh+ZUfzw6mICrhFMrARgg2zXFQyao8oHM0WdrI3bc99j
Qz1QBcfN8ncXx62QxDrX7eg2derE3h4cU48obV9sGWc4gsJuntmV7Bgpjc5VinRFTpxF42Qy3g67
4831zsf0Ojt8iIcgoOLWOVUcnhFk9V5vkp3QetG52LSOD7N2b1hBazA0yWBIj8368RJXLz8w6cOW
/cWr6Nd75wD2WJLeDeuxN+IHPmB/9NKswBHehLQ5MpUermheUBf3s8ikjIsMF5pzuzq7f82Rpx7P
RiRc+6zoO9W2klrIFPeacVZbrlxCZTIkI4Q/R3p0WbbHcqPbMLFVxfG2VAiAGvpMn1Y+yh3NOayj
Ob/9LrpF5f+UaYGTvlBLVQPQqo01b5dV6UZf4/Jgde99S6MnzxKQcgvP7T+D1D/j1qHscBgOF/FF
D9LNJbmp6x0kygrjliyyHq0LNGlhpX9Fg8CCMftxvIhlo6pwE45TGS4KvfqeS7XXWgp455M5fsut
qWQNI7+3qJ0yia8shzO45UQAuEJpFF6gRC0JCp+EsOyd/p3sJI1AJ62qh9CmbwMEbHg1NGJ3CiOn
NgxBajvZyuvge9odoNDv6mtEKxL667hklFIvyRPJXMhcbeRCR2WcaKFs26KI0rT0PlqINjQExCyg
krvqbBprDuUh063vVu5bWfaxb4AYbcsdp+I6si06XCqS/X5oySPIIxWL4JoWuU+tSYqu5bfDfn0j
E+rGWa3TI3lkDQhwhdWsvRozmTbxPy3V4Pip5129b6hAcU1fJA3nzj9oZUDb7muBpDBuqIt0BoJ+
d259exVH0hBtubfax5FQS1NflxMWLrT1/G3lxEhrIAyKQYTabUgKBvka9clS3xKVBmhLZNW4ONp7
dD6qjPV4NZZpNS+8aTtnkdW3Q7vIrLrAtbq2kfnmB3y4X0DSKPeS1kdgdOActJlzZ33gB8l0hmSg
YUkJ7o+B/HLHatO0uSyzsYfGBQscEHtSRbcMUJxXGdXLbFP4W1jVjxRD3DGf/morWpwlh8ynJfke
ZJ/fx4CJDuJGFB9z74+fKtMZYCZzVgGNI+DLX1wKp7QgEpm6ukp+qrnPS5f+cNaci2gfGDAhBKWC
QpDhc7E1YDPQiltpzTpi8Pv0TPbV/aW2/q2Ixqle8B2aKr7t7oqg3TDALEdleN2OSypNpeW/GDTg
AkBP2v/4+TN8imVf6aDk45O1xe5J3duMj5Q83Nu8C1X8VJzthuy1WSdNpZfrxcFJ9+S8pke/pVfs
eKRRjFAY2vze7eS6bS+LWje3JY8EM2rBArKJeFFd9Bwk5RWYEGpQ9/9z7wTOjLiSx6lWY6u6oMVR
ili9iHNcIuEfM3chNOt2Se7OgP4E8uxNOpC4WKSTPPlgDRNm5q/BUEMqtjTh2oLYff3B7ZkGuAsc
6eUQtToDZnT4dFfisqtVvp4IYnntfjY1Ag4UMJ+puUW6d8FjdhAwsHlrtHAkniOjm3vm/90QVOHS
D+7YL4Wwu9AJH9N7Gor4noFIMUg3A0Mz9higRzKaHqqNZaD8hOK6tKryevoNjSmaKNy5fYRkIHBx
gHqYxTVLkQ3Jb6zaSZ7E2tx/knwHwP/kEjF4SLLm0BjlRnqhyvW9xWfp8XfsQnQsORXeNPDhbP4Y
KkXLhgxilixkQ8ZPViMzQatmiYKy4N/1qiUqVZwGay2m6CCGhyUcRrA42EtAAFWxsgtuiv528ZRe
s141uM1RmMudnAWgCN785yqpiC1RMnF0L513or2OkTjWX0ocg2RHUlMKJhLWAw6dO+kYlMD/0/gu
UaaRlJEexQRnHvA6YEWtytA6TYJqYs3KY1cTr0xtHBNWej/XbXTaKoGtQRTYA5sAIbiQ0DfwRfKz
kUlmJDRC/BB2Fuk+HLCFauO0POygYGx1Ms7XEqsh0pLdM17U3I2DXRijpQiZNboOt7JVFHbvWrt6
a/pT7hXzjqVMUKfSDDjRu7eROmv1TppYn3kh6l7RSoB+fWffp1/MIDcVKp0HKgNK5lV60z6i3Mws
u8YONUFbJWcAhi0RN1TQ7BTnrw7HclNrch2Bee8zKVpWwHRaNcJ2FMpzxhW3/fsZxIZ4/KZC4CYR
hBJRXEeGtEXtaNZGEB4gK/Y5mkcrvpQxxaHDli2/P6Z+AIHrNqoEJPGw1lf/nFcbTDmcgLqI0xS2
PssbECVRHDsCMp+9Hnm9EduGm3SpPI4zDKtLAYwV16qbjqHyMFXpFMe7uQPKcChmIsasI2q3/FcS
wpPBW/NgcSKIQ9AAP2dvBQ44obglidXn3mlHuZVCn31VgUzr7Y+qCGzu90iRLkiij2ccEyGOpREJ
Z+kZhmaKL8dqqCly01XuEY3WtZuoUaIoe03/hpQJbkSi0nRxwaO5TtlCa57oLEQdjrW51Sml8jkM
sj1NWVuc0WMUGPu9MJjA3AkTwGQUabrpIdoi0dYYjGfWWfMnPdgxb/Lyqb4u8CoBvJfXqtJCK2q/
YB5J/ZQ7hpCMEIqNhTwmZksrF5DJxyF3av+mX8yWJztLdUlsU2fyQEzODDuMD1WMdN3COs/s1QbW
nAiN2in03AAjTrIPJYp9xb3QphwmoBauOe+n9KZ0Bnp6yV4uOQKLgcnp00GS4CG2XBZqMzAXUmwi
/BULiIL2epXbX7dbvkkGDFEPskPoH6f0Tr+4RlDxm8mvjvEpfLqkIqIhJ1+kVV/7WhQ5++JaCqI4
BFCV3YAv34xECl1NtRLlb2vawdQL5UYZf3RJF0B1i/DJigRyr0QktXw4ouyQNcr7MFGJj3wb9LsA
HHUMcvNVINNKiluEMQnLFbSTOnt77n3rWqTTg09DaUniWC4FBrqEqqRAPV1q4W7wOrXJHuXHb7LV
7lAZc6IA2L/37qepGdueLEHCBfrfSs4S2hPADz18sJ4fStz93McTqw9UvjIA3NSb/TN7kOjX/Nqs
TJkBt+bWor+Ds0ZdW0UGp97nYkrSEeL9dMS+KnDomJSQfeh77UrCpD3AtfKYpHqbFI4Wew3VbjEj
leKD7MPuqPhkjxoRnqvoX5U7SOP/FbAjoi+ssGvvs2aUlti/l2ZViu5IIW7ri4mlQAX3U7aQZ3N8
TIupbKvlwmUoQ44Pc0LUkjQzvrCG3NZ5n6tOQu6SZnTyRvrw+OUsInIc78VotNn9YrTDkJQ89BEE
4sdo1f+HUzZEuP6s5D9vDsZU5SIjqWLjvOzeONQAxINEcRwXT7kJhVEtBElNyVbA1oibWj7rTaZA
W/2X8DxWVtEEtMzj+CzrbYFZbAMJpX75m1zOFf7BScO8uMUl0Ou5jEoLIIyKWOfAqxX08S7Pmfzl
hrRK8k9jQXtZR9cqT53uk4uVDMcTWFL1t6+ZuYE2/nfXl7zHtYqYLFBShPQWrJVVx0r5ztqzrT5i
DZjPYhazv/I9qeYG2LOcQEULvwbYTyqmxp09FHofZ5/bukuRY+YrINelrdAiuiwGg8H1EDvXCe5l
NNfvrDt+vxFKIZs0sU7qxiotl+CDZztklsC8aayOXZmC1Dxn9JIixXRIsIYlqUVCg8kFpOY+8mhH
FuR2PKzyI7AjxFThlj5LLBiHEe6DfU+X0pJg/3RCh1mnpseGyeFRLH4vpqB8a9S2vD6gBJl0jl4/
4mttLR3VftlI3qXSju9FLVX/whcq6zErma6qIHRyxjGjA5p6CFpMMby0wlXNZplwzYnkZrzBZOOQ
6OfRqLzmhq0p17HSplB56LG5qjyfwZ8j3d7i6OKYitKHI9j9k2yR8hlt+f53mMdmhnR0FFgstO5s
ZxcuOtKw3t+ld/HptzfO9/xEYcL540CtVfrjPvHTNDQEVSBKOJHxQLnWDJ8lykKOW/1POFPqYHWs
Yo/+UVKGlacex5YGtkAtDU9E9QfelPh5GZ9rNNwnUoi/LNhvsc3JyhN3AgnkM/iuOEOds0/bJ4K5
YEd/ka3zvRPAsKfHi/i3szbUEAwCxUT/wzDugegHw9Kx4vmrbcpTiC0pUyTIty0xXdCNmFDdH8w2
gycEwt3iCJyU1pcyY6waYFYDn01+ZYtxauSaCR9fJq2ECnDPTHTSZJuBPoBoli/KZ343jrq2rkiN
uasi16EiAZmg4YgWY+BLYeoYd8PChzFdSkrp+xmPdzQEp8uQZQUf9tcsOau225/b1T3jfgsa9Gbq
+W0sQdQv7D+895zKtblU38WNg4idLWcP3Mu7wqzUHxGxwxkO8GFQpmjsnVqAJaU7LNnizIZGPzcV
lF5LCTFLkHjjNsWCTiuHx7J/sOr3zJ6s3dKMFoQ/jahzZzIu59d/YP6/+xLEkJTDIZhDmVxYtkYH
NJNkSa3jchrKms6J3JQwCqewFr6WhvQ4VbeGRV5UczPokGr3gNlrQoI2NcKrSLpEvB7jEx5UUCHF
asaS03+CSGqAM6zAh7x4nTfhB0eIGMhDVKS8vPL0EVkSuXBExgGFvAhQgMhNmIFSM61LDECu1VFW
M2xjfYnhrD+dv43RbHaXkzJC2fAfMjJUNROmkRZ06kzTOg8bmJWLps1hDaWTfNvoOWnfsMeiBfHw
T2vLhVMySKALmybvCvPDt0Vh85QXr80z/sfcVw/oyd4W7yV7gNcR8gLK9nvoiZiFb/chAGH0/LHN
yw7I2ayn5mx2J2nW8rmv3wg9uxs6PFobPtBHHP79QriN5Jimwh9szPsHdRq1CKvBk7HU1q/imvB9
EzO5VI3Uga+XlTOQByVJtEEPcFSgEZukTIV2i8YSSWHJ49FG6d9rJp9Llyc/8RFWuEV4YbWgPx9M
g6b01edD2P6U4uAq7W55fksufCWOMllCqm9hqwJ28g2pnaWsHMpzRU7HMFhdh3cWkIlfi1pXYpSB
SGcAMrvNFmdGkEnvf7Ic2xwOdaGL/h/Jiys7voF7NBgbmKi2FJ24IUFk5IJC4eOVP5ECzFqd5o//
wKlfmS9l5iSVO1uM5bThA/YYwQTlWZKNzVAufWCZ7Gez1lzQUkiMa1duUJFvJwQLbFCX7nIDxT86
r3pmOc6EYWACiBB4XMLVoCJnXXQe3EElwaXtUtO2sOXXmpZJ65x63x4tq3d4UmRA3nEpCvaKfaV3
a4yIEnPWxn9af6LqGlVKsjtVX7cejzKq9Eo696Nc5L0Nyc+E7SMfDoocLqU62xP5PDfNnW9haQME
BK1hQLXL6IOgPVWASslD9MOvj4rAWWWDoIt0vePAO9fg7eFu0tBqxnToDBcUcpWiQBIH1GT6nQI+
kYxdwSeamhOi8Pda/GwW5BwVOooRT5/UoyseTSnFWDyV96QNuCtef62C2drz6OiVwYiS2zuRKiI+
vKV1N0ybq1T73bmtR7U+Xqmx4OvGJm1AbECTK9uhFH1msj7uyrJf8ghwacToPExqQ3hy4+MITlnI
2q3LN5LPkmnNfKvRuqLNOWHCxJmUK2eMMZp6JugjWMCrN0Nsj7O8jXU9so+XrOpEZg4T1P9qXRfX
fHpCIwHcnVQbRlljn5ZJAAjNkNZP5C9PAPyxFYREZXcHhGnAKYwkr67+NoWRF7EumZ5e/Yn3Rz2C
CZn/EBbD0P4jpUTJwqCwYDQQQtdBv6pnFgNmk6IwCHt/hlBZiADq9rNzMYVJ9I4b/33g5US1EDKI
pa9WjX8kLGD4b3MvOATGEh+LoQ5PgOUSLwKoK28XPAGBJNsJcyvyf4dGImDQtA0AtE1BIFGken+F
0gSzaGs1JvI9kFS3bOwoSIuaK4QQ60cIH1W9IXQMv63zYg+FjpaSqopYhOOUjgvCwS57qJwrtsvk
4bDXW4ZBcYd6ajB61hsScbWdVZMwiq63wjE1HTJjzbs62aF/782Fpdul44u8ip/UdzWbZXqHp1gU
pI/GleQrh+SoXIEHv+NCKAyYT1NLW2tOJOqvIDc1EHszNb7xxhb4XddgIdPMK48kSQlgkLSRBuYT
aiy+IAO1StfZJ6gWcemGeJALZToPNb777WiOrejRBcN6QQBCKmhnT82WvlQWhf/MxlEgzJyzGbcQ
rg1bJziJ2RbhzSsjgZPlkqWp2qwWM3fpubAN1fz1Z0gYlyRQK6QkQXBcgdAzY3vOh4MlDtDjIAlY
0IuKJ9Yme9e16wE+gvosTMaHk2r+eCLw0QAxmoVzJLEeqJ/Ayx1ssZGx+K2DCGeeGcDy3eSDeCY0
fxdSUiIacublMsdWvnr7M7oEK8Ye2hWKQJC2mIKGL2mHjU23rYQalMeK/I1Yf2sTBJfAUO5bmc+e
lFlsW7ELaxTftz7kuUxu33VnfeH590rNyPID4KBhvYVOYieycFssXjBN95HJnRUpfhioeXW7WwCY
VXEWJP4hrE6zHCP8OCtC9/b4akqpYLLFVCZXz8XO8rHHV+bFIsG7AHsYzPntP3npb+NhVjc8Sfl2
ej8PAA8Fo0a8afYGee/sJpyTC4JSxRgiZcu+S/Mpb9AYiO7CNerdFWLvqDJYqm8DiC7YfvsIA+kn
ewKPl5wozPg3Ey2szCZyMIf9hxkUenPZWwWNs3sSSi+EaGexuWtrmYHD3lvN57hQf3Uhl080HN0x
21mhxAHIqIDBT7I0AS9OBC4HPVxhPTY8BFT3sp2CtMdkkFGLxidJAEia9Hw3xSTxrPqKUfJe1raL
qXP/SzJRs2yXtEnSgwcSa8ISHLwgbWEQOJPu5KmeVwcd8Qq4if9ZeiRQXG2eDbqRCc7+amz3FKfz
XJaZ0vVseySm5Bd2IXDbRoUFfojjYclZgqc+XHeesNhfSiPT01gxiSt9uboLtsRiRNttcdhxAb8/
7QgWIAZMn+w7nhJ604Y2d83GI7rDvl2M4riqcRL0uMTHEMc19lBeqko07PUEeUV+uL2Dcbjf5BCE
rNMJ8JAAWR+HKsJQFgUMeNmk0JKR6RvQfyH/h3FBXVvo4xzQFeg8yHPyvoPk+DIuT+gveyls+yXF
VJwPNKajGVCEQ+sCbMFrrJHYoTS92wnFqcDtyMwPLzNqmjLUpPRt4uDZ+hK9E0kgFQdLMbzI2aem
alHS2lj3Fp5+O+vuFGnA2mHAwWMIva4LmkdqwCAcaaunrtYGVw/y5Rw8DSIIDiECizV57Fm4EdCj
P3wLyvCfvCkKVKEjwYWI4/Fh88BT8a6+ON2BSWJZvW7fAeVXXRJXrFlRPxheqap3oGJrCm/TKmiP
i9C51wdvJIhj2iwoIBXNJkbGo9EyzTg48KRU1UxknRPdLBuWFZk2EIX+ygg5XImPmJzmsJpDulGr
OR5UEz88r6IKmPdvQXLBSNKfuAxEZdI+mliqCo3z5W5vX2EkBKd+LRL12saByPKniYEm1KojDS/Z
+Fcg/Us/NY7rr88cl8096lRVVB8fZeTkeknjpFudH7OqnZ3KyMQ028pQWCvRRnfiqRViOOIBVmzk
fkaQ9sQY4fJnrB7ZTu61vGm8oq083PtaHlA+h5LMEzUZyuyCBKryaEuntv3pWkRW4NZOpbP0nu9x
TjCTiapGGOAYUVJpWzeiI6PmOiAWxpnY7v6qCLdqiQHTFtdQ9xvaw2GF+EtVCje8eOdJtUASCWzA
sAgKUyGfY2L2ixyyhR9B/KrMw+ENcrFwXKjwUFy0TOIUWJWu9PdYMldRQi3qrdzUzhTkAEGlPolQ
9Usbj3Nxd+RCybwI6Jj24cMsihNvebjq07DMV1h29HanXeDx+M9r9OFJKcp6DBfpMiTmMj7uB1M6
JTIkSEBlYH9QjGERsVgE0+6kvs4Lx0Bbf4jAMspRXbN9FyCQahXdiPLEJoVLPVLeA+U+EYquzkjJ
Y4C/8agF8adoxS45rOl1E1dhxZKks/a0661G8l9757P0rWU1xt/Dl4iC93F3SabwhK9S0+ZCwYFt
MFUy2AYIxRNBSO6jFZLcV4wAeOs8uu3jqqaTbw3eq283tdVurt/a0ySw7iXJcSiKxYzMJfFlQNrO
j6X5JiWMGdANGh8aZaJ+zB/k9A6EGlP7OPes2w5pC1DUbxFU/G8JEqEnkj9N1Y34I3v5IQxdF8MN
VNAxQv7uBKHS9oNY9vL2+KVkApRC9meKvGsyqvXCu5GcsR7mFvTh/0f7pZoeGAON1q9JER/sbzM9
/oJtdW9jKbPdN/HrvvhtEQCPFxMw11tcN0Jzub3K7v5qw2hknUrxpehjZ5ryeRQjU6nc5M4fDhdL
H/VSBWuhVpekTsqWlhh8KPd+arVkwD5mqaFSNJvLaWGJHIVsx2u90+FU6JUbYmpIHwZr7muBMwP+
YcNk+pedPqFEUVUu8f9dYhYluNsepAtTpBlKBSnJECI+PnYb1NrVau+hxDErtltIVwNYBpa+MoF5
JrU4mP3+7WfUQBsMB4m613TqwDP0LXG47v2XoaU2v0vc8WWiUcJsRyU/5VRYClfgCnbEMeBUDA7F
1PurgC6if3GO4jTULhpOWRfFznY13a25PvR1D1pEZPugVlX3G2LbNgwC8aPIdhRr/8gXLaK8+Kjj
sOdL8XIpxf4gNVtvLgY880ew5jDbrZx7WplZATjefcBQC9UwEOBGamCZM7UUInhheSGbE+EJaLfb
lDOxi/lVuzwY1i/eVubgl5aiFvclet5/vGetkfiOFbxyEEZv58wKRmQUYdXbSJxE/bpFNiliosMD
h+OfdkZ63x+j9NS1/+7m5JjLiOKTZ89z6g/1DUeMMWzEuZVsvn02dpKa59+ZmkcPlY3KNv94Buvh
T3R2ODmGigslDa+RpRaoaDTtn93sJlxsfUYQBiwTyCYMNC29VnaQ9G6CBMD3lljChx28gaqUFigz
vWJuLVcxXgA3d6uhYTjdO0wakx9/eqLwIG+nekI0H5Mtdh4wG4MtaS52p1oaSUbC8Gx2mxWO/mqp
oDsO4TK2xkzbUl2rZhMsQihSBTGWk8U2QrKD+xy6QfX2YirYkKVSjSUvA1MpnLuWO4/XaQSoYlOS
E2y/Xz8PWnhUe+FrfTiP5fZ4+C2KtmnghYAqcYa8mu83W5KBhRi6loHpgnAoZPqvgEcJc0LdP4PI
X44L3p38GLSkorK5leY58at/j+5FD8UwmYh+xsT469+5ul6Wi2j4Twluv8cqUkFvLzvvFfhl1G1h
Q97iVfBHorDcwvdw6dmQWoqZw/BijF2eA4d6QfVfhQxCs5RAvFztz/EqIqPTdbq+BWKjUTfQKJkR
T4ufp6gh6u3A3AEe9cAeX0Q/0Vp2X5L/MVCr6F1LhoQtfgi3YBxUKiPb4qaMyGfINT6aEUe+k28T
dLNeZJxqYXs0ZCY5TMXabgduFCaZ6KdiTCyWU+I9MgcvzoyrCbG8IiwZ0PxsEQYEQPkiacbsoiAX
imwrpF+860UFS7Jib0COPwYZ3CUbbD0oRxXdXkqBti5+PLzpEBqbI/2VQF2zUJ7QnOkergt0ZbJa
pqSJW0StlReIdDKbM+Kr8LJbWElUeSoZaAXd8FJvo5I+zYS/bvZENbpQvV5/stgOa4G3iV+rSH7z
dMiHr6HYPhlNFta2ax1lMIYTXhSLVf+LSxWUizTJqXt3YsdnRGtmx/Pqi+5g9YDBpjlYowmibWTn
AmfSAnoFbJ5iXC1CmtS26fx8U8yzsokafv+q5rBSWah0LzWdskoVS/PbzBZdOwurAFw6DEqJI7SH
xxO1qjQ3Wobf1DTzMGjIj/nXaQU6FcV4fxxsjw2q9D8GJdLJ75wK4tLq08sSwhG0tMvZp2MvD8kU
sYN6pxJMggydr+IH8NMTmP3VaSnW3EyYwDY1HDzzalVwW5sxyOIBO+U/U3jN1ETqfStiZXzXj+A2
6LhpYq4nM0Qikapl0NIew1nbsYy9uwXvI5GVXcPPNzh7+ZUVQ5foATMQH9ALmsm9S1OFmrJdEuY8
2dxn1jU4uXOb8ySkuKxjmaTJqr9G0jO4GlwaavXcsfw66HY4amaC4KWSBOfbNMIgoUgQvVZH7tIa
K7L/UhG2/o8kWxpoE1olXyjS9wta6zr83GjsomceAfKSStzNPSq1DE3DgYOYSTr+3de+Vv+ZauTE
z4XryubeDZqlXilsanEGzrZPhGkgCEgliw6ri41lqj+JjhDXjyjos+7fWvJ0kohOgzUiYxiBUr6l
ndgD8j+saokI9/t1FEAHVV0rq9ONQP4V3k0woGBseRTKA3GzGY9MakhNgd0oUSXkvVDgNW7NXY8k
HKri344XsoOq49mfraUWGk1oPPLg820xu1TJSSLhx0cgsqn1pyXf7J3E3Bg+uGytmwSQouvP53KD
AjZzQN8k4zHHoGYXdSebkgc4YpnZLPOuYEwF8n5nuGEfXcYHK/148QodaFC0sGq89NyXrir2i8eT
TayOH8QeKFsS9dJvAeYU+5dcvwmVKqwcxTgonISJRyYOK4DK76TGbYCYgg6pxeamUcclvjnQng+j
0Z8a1So0hXU0spPoXVoioffZzprZmMh0/+GygBhtR/iDjcLd3Pth4+0Uobet4chGKDi52jhlvyZk
rJDGGhCl7qHNqMsOVllmbbI7MfAAbopv9El7bK1JM5Bu3QkPovxFI60ELU9fV50tyX41vl5CJjDD
m08tFKFZXWHt+u44a6ed3lSdRyfZVjQrQOIhRdHRLwvOxQBe9PJ2msNMbfrL2Ia6cAH+gwgoepH8
pGYSqcFbhp9j4YYVqDYMs/LeLOdEwQoB5epnSibHP9SUwC70f06UNP/xxd0qmLP7LOUBz8oMTxS+
JeZ9Nbu4MHsRhkaynlGaSHQB54SZtuYmtUzo3Ra5R7E07GeUWvEhP44lByaDL5I0k87zo/CH2AZL
TmZahwqoEBpS4OC4I3Xwh0on1BgQBpnuKC+kyNHaBCo/3+9RDOxwD1MNId5uMx53pH7JT5XZirk9
aNWGTmdsOM9fseriQ5RVykBqb5homYrEHYBcLJ5/fDM1OeIMhTTsr1ll8eCPFmJjPwERR2p5zLb/
V7UlE1kYdDHWIxaHSL1ht09Zo44iVMUxAUbLF7UneHCTTvk0Rq1MlzHN4lZjjqMNSaHEv6JvtMvv
8zIbqX/MhDniRin8Zklav08Ju0FNDkpvXCsoagD0gjSewgKiLSRuL7unKpsdg8/jLYMF5fC2Kfzp
P9hV9jiBETCIQhtA1nf2ts6msxVZk8jpvrXugMLpBLf8MZDbc3bYGcXq6Fi7ny2LAyKr+WFliHzy
jwsO9L2wDvhxCevs/oayvV7d/OS+VDUIlRk3AZCOblNq1FlqYTqi3CwPZe3zFZL2CzQr77ydEkmd
bAI/2zf/cqtyoVq/IZgq/yTtfx3QZlXauD2yZIkL67foc2/DiOT/Pv9oio58Rk+gqU1392XyahoS
W0ivNuLScAU6C3jO6wKEDzD0jz7yeWnINyUAZiaTrtR0JgHWZLEr9As2rnDe29s0DgOlgiTTviEq
RpKhqstEGRmZZgWo3MGdVppdE/d60JI4tfzRmQ1lLRn7im1Gt+3XYPh9Tg2aIir20qXMXvRJU5/p
oS7alY7YEEowVSHzyj9czqWAlPWQoMI4fbLn9RDlV2yjGPWHIYAl371TY2ZCPsyKItS0GEZi4krH
v8rFxkq/RqNPx6dd9Ja2ObXezwZ0IL37ALKW1Idd5ZA+eIBupozS88QG10vt/PwQevHPfChVF1bH
eZ3tPS4CcfD0WAgkTbCNOq0Z6yIK+EoUx26Kiy9ht6uF4X8iHTb/uCl4U1ZQrn/O1SQn0kgqmgqA
cCvJxD7yg5n2rEaOEBm013n0gAPjl+AyU89e4+lgOjGliarxUsErsGob3QgQD2piZx3TBAbh/Iq9
4B5/XndxQptyD1EbM4DgHwgD/jojLVZdyl1k70oqUNFyb1xQMIybuFcgKAYrBBW6GipcLYaYJSNc
5iXBngdEzHyq+Sna4XeM1SyNz3uadmdOXlIwT9+VFDoanr+x0GkMnZA9ed1Lgw44+IAq+jHYmp0y
yjRIYfsvXS/fM/Ajr13G5L+6cppWHHu3SIwKc0EsDrNQy4NXOr3MeLv1OJGNwt/TzimQXCEXVW3z
2ENxiL+PDB4f1DA0wf2l9uEr+g/W3lfD9MEdzxF6EzFb8SxfNLNqvFrWDd+JUPmHi1vbaBJePbdg
evPsOVQ/lOlsswpTygUW5q8rzniVcjfsS7wL+hKmmfacNpiSictNSCsJH4CZ2PD4PB7EqJ/PNozp
GqY11ZjNyzzEDRgz9WNqgRNwH+J/ilKl0Yw+lQh2H1uGsWSAdVz0CajCTQLxddGUUmxOujcj7j9f
mOOj0tpgxFWNV7qU77zIfg6Zdk5+pFic0LDKTlwpc38VmVyl5Cn5OC7GVyQ7nGMQC57KWblyPN8d
2uEd2G9jDaf9sCugs5osUhNElNTbK7ItOY/O5iTWLEaY62IzNkFehikJU4VRM9TBXskl4Ak581E/
0rvboA2TZYZp6duxOLCnji3F1e3TI30E2GFFJRldUsS8HPsAB4cpgBMd6oWFfa9G8vGDxLWQKfD2
6dfWw6SEQYNmyc6ocsT5BQ1vgbjqvyocifqm2FhsCKs5QL+51J/FFyRe509BpcUDPjG+FbsS2Tlx
4YGFRFARngQpyOZCErfA7oBWdkMbo8+qfQ6J/PeH62NcxbQVXRc49ynD6T59Zu3fCfrlio9AMx6M
mM8dJLD2TWGQq878dIMihIMvl4lNMjxBglcZ0Q1aRh01n7SnsUi01X05lwUF8TJRgTj98Mq4SF65
78H+YwwfY5NVsmIjE7EE1GjtkWc4BB7sGyGtfeQEEJ35KfkzFm7UooKIhgyaL8LluZXahil1ZM/G
cRNQ7+d5bA4KQiabRQ1xAClG6Sg65uZkGXko9D1qTmb5YP0iu/ZlOfpVshTuy4ABf6PpC9q3MpYg
iQO39bS+0HBICSltwCIQzPmSZOKG45D/axidSW5gzzJBk6sU6cuwnySIPuv5s3WYau2p9VbAJZV2
S8ZFnJimfMfa6KDgydVIZLpeEGIT+/ht0kj1US0znNEgyy//ZgvrF8OxKbzUVrDSNFXyRfsUpQ4X
6KT8QVID4ALETNNswb0EyYIHzX0hjEdgpWZh870luK1CK+LrxZE3tWJJC2MESNqheP0tBaYBNkWR
vwnwWsLJLrP5ktdw4psDjXJzxp9q92LWfAg13+mePbl/tFi/SUhyV7clRKJyR0lBj+e75FiF8tgG
XXkLxwKFrGVFQMyBfgSyNJVePuQE1BAFVDMaiS0cX0MZ4W3XmUCBLEAGByBPqju2KQudvcKtwnFW
3qhdJq/gLwa6GbsmFjTQR/9quNmyriyfC5LhbzlfRkNRTjBJBUE5tKK+6oB8wQPcJOv4GFrci52r
SW/U/+GFtlRVcZIB5HRwSbL+ZRfZyJ4cXzSD0T475hsjVARhO2YBEHl0IkdlD6XrIOx+LeeuToF5
3fYGlhRqDM57t5cW4FLdZ7yIKRaisA9ijufzsEpEmntE5luztd6wJNdjCnuO45ulTa+EVt1PoC3y
mEKy2fUs35v0Re2M6JNB7s3TNKj7dGK/NpLLdRh4ocqW4mDTPCqYgx3V0/hqRKElhX0YLdjNchE1
xWprMf1yO+ElPDAzuzp1h9yBSfnGIxCyL97uSCU6wxgrp+ksrfFEphNNfRJLEOEbGQk51cEbhRkA
5YUTJjlAhLcItkHo/WHzmR7td9zATESxY4IK/ZdynBFrxWtaG2Gx1kGFqC0LkArULxhzQgi6ak4J
n/HIjSx+aSSh/5tluP+ivunTj/5OE2QlHf4PRfaKBJPWd8fMPpge5ayW6rqGW0k8/fOQGLo0BXW3
gsNTiNtZEmUezKjHi8V5bJKGZcdPAkiffgQJuHQ6IRPR9661bt2kziE1e84va9wA1NiShfcqaKeB
FW10Fh0htirxw8AIGjQJOcW7GfNtVHAOX0Z6FvgmTapIsqCdtuHAvXCD7CsVrZ6yxBZyWM5dsA/Z
WfexZQZeLFocgTr0lQkd7J9RtdjHZmrY1MmR/2AhIvwyqzcX7eUutoUOoFe57UB8Aohu3I0b7u9V
K8D+aXpCOboB7e3X1xVYDxfmlLejso+Hv75emZe9TSvsSMmXrULdqUu8qDV5ZpZkiJf/HXWyHo6X
Gz7OdzpNc8a9e0IDE/SN6IXTX0s/2IkYkbST5ZWISXxeeVEsK7jdASn7aN1h8ltUvvkAjzaO3d2Y
WB4EXwdokMaAiRcno5lu32lfGFN8sgvQpmoCBefs4KX6U5YOpuAwQ92N2f2WS+YfO3RKqKtHWvrO
04qSevWTNWfLnqRfu8KrpS/CZkdEQNHLa4eF4pexof4F9DrBvRa4nMAfLzK2ol2VCRBvyYwZJ2ka
weA0m8dSKWqi4YlE53WQysX4S440KLIoDCo+kYEaayeblH8ZzbXP1Pq4TgomnO7xJnAuklGV9ieB
VW7OU8SCdbVBCrAJtzo5ekJBBF8886xaPnJRyR/TWulVc4R67YQi9+90qKucIx1pyDhhZrNGoJ7z
wZYnwPV6HTrMJwNzlNIqA/HbSSYb/AixoaoG2KswBBWkctd7u0PbJ2u0950hrEBhzk9iWUfLDjhk
dDDccENYWy0rUBNgtQbo7skU6zQTnpFAfApZs9dEFk8137m2x9mqfwjLKgTmnCy/X/6Hq4ikvarq
+iFgcOaYTQjB9/eoxv432ilGTZwvTvzqirie6VIndsKasmHlwHW75hLGbewiGPl9PyQRXIJNjMiO
YmR5l/+cWYX1iyd23+dM/ujNUs9endJG1wBMZOctGxoLBIRqmE13a6LhBJfZ3A2hcZ1/fgXIxLBj
8j0PlQd/AHjj+h2G+qO/UdygzsYoE5m5zkCFgdMZzXIBxxZR12YVwok+jjKCtFhYGswjA1hm187N
htrhqx1W0dGAQnggYek2uCqKf4dckCEgKESSjgHGZYnoN+nbbFbh273odFFWVG0lBfJVrsnp/beW
yf++1F/BGUU3DsdwPRetlpTsdbwNcfbKoqpGh+QGbkCU3jPvviuMV1qg2cIvdyfY3x/P0dIPulEk
nrGU8BedqC0Jnwwt91J+px6L61AqO8/tZZECCGyumIYtlLEN8HqNTUknfqGIhIcOnD7nAarKhKnv
DgeURIaLTsD0URY/b6i/COoA6pC8qtG024hKPoG1w5ozZlk4NDrHzxPjhEe2A9ndANOfUK4bN7Zj
BcIgql82v5P8D6nsqlnQ2wkmPVWT3w3jfLDcEnCstLcj7KwSXZQbgPNsgQ8jiVQfU6VKktOqLLre
D7vlYayj+c9yA/XM4irwRhhwA/kqMh6M/IEKf3S2CE+t6/790se/cL9KMJ8TXnLsf5jPxvFxc7pp
vszsX58efx//gw5jaDVAeSQNWHrBmrzaJRC4dS34Ba2Y0Hb0o5es+mJcdZoKizLLl/nOCdAmn7SS
+gTmRGlj+ncnnUlGtriLhTwGOvDpjsZePC/+f+uV22dp+BSx6uaZzcEl+D1KLT7y7YVyoIn9hYqu
PSm4BLI5Fv1DWfw7MtPSQ1JmSKzbtt3IaGr3IWMMnJsFGDgd5oDhXGHIaNkrhDzsJQcRztH85QQF
M0q18xMtm/Fx3qhAKz5YKWbIpD52ycI7tITHh0AGzWkeeU9mumd7azK3PbsWrZzwOGaqI9dbIO4J
O+jIwNO0f+Q8Rr2/aN0lMQn5AsGNboQ6jHJBQqEKkz/LXC8YUw6vzwjOuSPwuE+0TrELjQCDmHNd
84NjP9skOa98zmVe/NrJGgSRCLOiYzJPx4Gt/ZiyJTAOF/axxiqYbUuNdGd76cJiDYWnYvPhZdhK
tfI9DeDdZbFMmT1JqDF1sUh74hKbFE1wnF13XJTQfWwMgdlYY9MlEcYkBToCDuV8kGU8o/feaZ09
fB3D4pYbB9WXTMFkZJK1E+71n0Kls5kLBO1pUrUxWD7J+BC0NenNktCVdNKLY591xcQK/oMGtDHi
aNZYVsomuMp6rxNTJkxErJJuuN/3jpd7rL6l1qxsGb/SiQFu4B/H6nJOzhpDBODxogHxTXihif7T
wSWzyvb33Rpmh9TnghNo/v3vFySjjwV7KVBYZcmHch8dqckI92bejKYHxAhptBEpxmPflHjUDuF4
IPmZYcxl+6o6SKP7OBfmuItvo/2qFHIrHDtLq1dioIpI3HaHa0gTtHtr18Ftq9Dlem+vbNAcrkyu
3B9Fjj6j4z0OcrEQsYiKxaGkY09QWbpTbSEnz8cmAZplv1xyPV+YlTHG9PKh3bLHTlU3+jODHV4e
FFOnaZrlwlNZcML2soMTiYQt0NJUr39D5GbR5iyUI2PCf8GpjUoMGd2IM6/2Gfr95ABaKhSwngzg
4iR6tOmGV/Yxp2LF3Zq457fEaCFeMq7bTh9TACTTkAe11ijlF12qFW6k18A9Ug2p9iGDrw8vi1Lx
KQ706CtVRRT5ncQuG3EYwX4URGlO1/fwLDUeegZvA0/LAfAApdvG1tTCm7J7A94w1gPOLzHAl/7f
JbJXgv4BTD8SN3NFg2wqU/0rxSRbAd5fXhxV/VGq9fDZKZFLgXRGIMEYVH5fLYQ571uPQVPFWhUP
j21zfbQgkl7v1jU8jPmlpb6x+IkrHhh6C337mvfilf8TSJAguZR3lim8Let24qdgKF8g0FUqb/gO
911iJG9Q2TPliPyAmr6hVwk32/UfweLY8tWY2Tthc9sg5adca4UcrWrig3RZzngP0eig3B8Bz1rc
44tTcbSE0tzptBJyMuP1yMnPYUuUhSgTZMBMVB14KjJarrcefuhNinGtZztOGV22gU4S0+cKJvpx
UOirHcc9Y+HVpXJvUoqHFCNAlC68d+D32sXD6Qi7w16Qo0/OCsV9I3Q2P+YxMI90z0MIk06ljTdq
Dk4+FK/WHVZb/iXeqAKVg2/5ieN+n0Q3pTeubSA7mu6ewO6Q8tk0XCfVrmvNuWIf2VwZ8ri/ErM0
Myss5B840mOWmbULGg4NbEsE1YkCYIVamH/z/tbfjtDNddmVVsTFybJf1dSXO9dzKN1AuxFWG3KA
UgFp8OtHyMPEzr7/lbdiuX11lom7sGrYnMN/vY/ncBwC5fF6e/Vh6hAXIY+1r3H91CU7qCZ4VjXN
AcZydSYcRIWmtC3f7p7BwtX89fVzrT0JiE6TWxch6JdfYRNOc3ek9JQlChXrqSVAA7o9AHLUs4QK
7kR/7d29LaQEDkL4aWOGutp49Zc1tbmVbYUjXjaCLJl5kE7y8TpKi78avcUcCfy8EU6BUW0USirQ
E8XYAc4xVHlUAHO1z0JK4VFEyfoIFuWof5tCmkBLZZRWm4F37mjkPuGSOGTMeHRKiHNX2ibQeIQ3
eZVOcncX/p/RacRHHWFgEP9+JznRKSCUH0WSM9Dlbi3UiAKjB/jSFcpYWTuK6/sszoUPkjPP9R02
nu7HOHvvAem21Y7y525AWpDeRFz0XdILnLO2y44ZK5Rxe+pDrbbSPSJwiB86KGnoui24rCvSO51B
T169FrIk2TspovvsMZ7lToxBK8BQqB4qZXVpam+wSX0m9R7Exj9Rq1yjsFivLyEWHTez/lm/MJ6Q
T9EZCaDtaUdbIiDDYqphqG4urUvG7egxY+U0AjCdqt6TO70tvxvWdmXXlW7LJqbZfUjkc5TylM1A
QQOfeTAN+q6qFy1sAKmYkylo64LMRRf/ypEPMj61zxVz9ti+0WsJPs/vrj/fWWJXbb6/nrRvspiW
lQdtiqKzk06PVUdgDs+bv8zmhxh9zbRpGVWWMfqcTspFZl6XyRK5+tFWvF9VHbKS7p1ggRIubJic
dMRJZx9TMSMaqlIOJyoFlUzwFCz9Wcax+V3i588pcNwDPvG1pEmcxntTtFfjk46pC6Io9ga4p+6q
7aG59DjbWdIPXDA3oYarzpIB0+DqkhtlaqVPsCOpkoqEiJ2f/3Kx2x55ECvm0R16oRwBAvmfxAPN
KGcq3SANOhlM14kASIyWCb/2EWDMOiE0d9mmDI5YysMHRdEGfRn2UE7BnkElhOXWQgt+IQeyzORR
XwmhfWi9GB95ME7qScKGflJuIqUN5U/WipT+simf6iGJFIkQMhNMhDhzd+h+M6h5peO65DGq3YcP
4zsiFleoCkSXaG6ztixXy1K0+WsR6LBCaGKTvkeWLluynqquPK+XB4UqBnPZkZPs80suVZgD2fyn
1rZqREF/9+TEqZxKMltVJZXzMm9RifVZlrE0jshMsVvxXQFxFJFC2oTSrpe9uOrdqjTlZGqdB+qc
l/jvSbrKZTHeDbQXaZ9wSxXsimZS+kvWS6KC8TUjYFrGnV2BbbT31dS5Jm+Fx9mS+RklaXGMF1GI
G9woWM779iAScMZIfaO6cQiD8yN6QId10v2B5C9icCT+jwPTx6ipxPF11+Fa3k1wv062Zc6reCTB
DmEHy5uOur/DUeW7Tagufr8QIWspefC4UGbM1fF+n3YfESgJ+QXVSwR9TwtPAh9z45TXZfWSJkC7
G25o+rfDjDmXYXyR4zYVkB/P8HLXYy0xt+yqUVswFu45UiecpfN9wf9eYfLK4EYR6WaLTacMGFSK
QK0qboSeIE3Lgcx5ElfA0K1K0fjklFG9yiuALHijJUxy/fS2qVCyR/FLt/jOjePW5Uk1YNa2Wzqd
u2O5J3i/vZHuJVGAu92THnW1eIZBPd81OgFzo4Jb53Ozk+szMOh+R1yCEWWVpa9/AU9QyILv22po
D7jiVK4/2MelyCdM899EQymoPH9hR6vZYgMafdjRIL2+995H1eee4FRc9xmamhRvdBFgS0BCu4xW
ia7KDkYhrIbOZL4X72kBZpsxQevvnPCKIwi8/60RSJgV9r7enIGiVxN9+nT5ynBO+Ay0EN90uWvJ
apABScA2uXlffCMuu05940crIGJqYAmJYA12vRP8i4GGPN+16qaYrEf9uqt2gGCpxMq5qrVvXogS
NP1qQfu68H5tBkvgnlToFmtCm3hbncVwsUgPCekwB6J++8SnQSwDbpK85Skm/Tli77OcRQV7eiv8
xXADpVOPqouqOniKTfkSmXkkNM3Jf6oJfzcSh/cq39Hg5kdVVjHrjG+M9jMk0LymMjeyvP/UAYoH
tbxnh+MqDtvueFFXjyATJck+k5V7rDyNcV/DsSXeWvGEXlA7mpj6J1k8GXDqpphQ9+LFAE1xebxC
vWtArEZn6ALLIf+dZzJjjxXQR732LGuPmmIcDLfOin/YUyQcdYDND7sj1yZbiz81YLg543uBeQNf
wtrfCx9OERiN4x6wejRJph405wKJeWV93JJpQZ3FloxhCl4SkJmK6EGiopMnbwkrSJwv6sXo8gQY
rYPDflBUP2/tFZShsTK/oMYkB7YCYhuclVJuw8UYMuvG07G2xBuaJOTL0cSHjVD157oHepk+qtbW
eGj/IQB8Dnq3DN143Xh/By961j1ZBFwZUxE1SFUwAbxkvWBVsBqI79DsjTRpwrT8ZLAm9KFLKvQQ
SnifISoRt8vJujpcSJA4l2nQec+2ISgckqOhuvNFgTOWBrIhl9azWrKESEMzUtfLd87gb9onW5P3
dkYwu5JBrNIFDlrjh2aLnV3mZrW36iaatruoKpfc+hJjijYKnO4laSBQ1tCV74pJPkolHv9q6Jws
RpLU/v8BkMbBFf5yOjl1gdMYZIxjBk5Cl2fQ0Wy5utDycy6yTRC91Q5eC1fsSm8OEDEWjHXwhLW6
amne1NidTQGrHVZMHZROQq9Mj+//b0RIx5Xe21Mxxu4h681jOTtm4DMeGWG8dpi3y8lEdGHz9MSH
KZxeERks/AjjmoWzUO2RU4xxV2PotchOFahTm9fFgHcHX4izDIFDyjESPa7WgRJI1IAaUZujz9Lg
iZpRMAZ5PBPhxnnp1sgPKAxs5mgVrcFmHfpJXaNWqNF6wxhi2XrpV7qVAvaAP5rXh+qj5g+nBDTP
G33wcSTlRIqRP2HJeFXrdD1YarW9I37Jj08pSkTuUgB9kc74OogZEV6fT4ntG2qO1XCqymuGsqcZ
x7tEJxWaWDxAsnsdjHGmIMFCqY9YNPTOTP6uzBeKUcFXnBsj6R3nqjeRlwV55dkpEu/0zKOUCIjh
oIEbv6TwM8ba/i7IlnuMfmLmGQZD7A2SLdCyRLm2xo8fy5RJaA5DWIhgubpj5eR54Y6bI205ZYOS
GDYwnlmnSznAI9X7bEPGKpyDpzeZHpVVN0AnSzmmwQzWzn4aFphMReBPAza44E+7ZvnKxheCbRVE
lmLrRwdRu65cK0ZkdnyxxfVvnw0QXv6NE3lMwROtoGzYEsxxMGa7ImiVlq30xj8BpaR68+xGcI4Z
/+hYnf2myYMkPs/2ebZIY3AhgAHXvP7U69OcoL1b2sbhgcQ5BiMtjotIqA/hDKV3Yk0z2eXr2iS5
cXOvQvWvFtq8MuqW4r2W3Pk/tV398sqxRo7tvA1K1iAGTYesQkLhT4VLvrgbWW9hZltLbQjWVck5
9LWxHEZ53hG1np6ZuB3IlHAcYYuss6GL3njewhDU6erwy2fWKm+VAD4ui2jkDpO5mFsjBQelpFMD
FaQy+hVeA5cUvtHBYjccs6XIoVcTGX2+3MmiHzuVAzsssTVha0stru3hyT4CCu3b62UZigMSWKt1
GTit8F8QQdQtNsgJMUmgwREjy0lUUUZJZ23FpRf9IEMdzbS5bhAPTjQAy67WdEpD4RQ6qvf80UZm
EqwsMo7sByymrp7Nfo930Dp9iLBPBWrnXmm3G9OBkgYK15zVG8qtD+Pp+DsVywWaaoilF3Lpr12j
D7clJOfschekUpDLGg+k5iKSHC7B0XmzG+4usoi+AGhYHFANcGDab3LJ/cIPASMofWyy+Uh0Xi7M
cPVNmsCwaXFmYrpNUdfn/Bx98P9kkAxhvJSUcsvM1FZzFr99BNs3Kw8HTsSPPvGpXCiHSkoVL3TK
AFGLHqu4ghyoRSUNCXKk4veAp7iOT8bJyAZlRTwvTdf0cyPz8ik5rROH1QKuRhrv8WmN759odO4v
3SisEPTmpP2pNtKNMtBTfVrAGxLrSIOdO2hWn0S2LFeE+q7+HkL1mr9BQTo9g3eh/WICIoE1y1qk
k0koN/Q0LqZBkK2Zg/6lEIsaTzrxxPyxrEjUs/NdhAxB5pi8X2eJ1Ou8xSCT6x2U9oETUihtqYnq
5H6Vp0OWpMvYNT/KjMcBUVasFTPTzWu0X8ZzbhmfIe0Hs5E6a6iRJ5yTlb/15oeqqdFZK6zW5BKX
GEEwTi8oyFO+TCoz+ks/uEYJvAJ+rXBXomHaI0pEL5RpB/MU3ZLGLSWfp6X1HgfzLXux4MpF51YA
3c0H/ZzwhSwBHXWSkM4NYKiFYtg3V9ef8HI+hLuYUPGmgsvd3CKWo3wU3W6M6p6PLI/tyuZjxxDM
I9eQxihgL8AGnyF2sX76HnVMTs0pg6c6kMuw/CeSBOkb92FjFXmzDC92QJVgJTrFwfCYjnwDxXm+
azEZuRfksW9goFL7oMztN1GiodgNEfdQDQQM//Y3/NP7SjE6e2Na5HFQmMlPihiFSvHw/fOx2yWw
wkfULxVklCWhSkv/DkS0DUrwSy80Fu4dMp8AWgMXEdbW5BYHEY30EjuIRmr3edWuSQL76hqFdqs7
pz+qyOSz9H88edMMDmnmIuxYp5cMXrC8Gbl7nYHnlnAGmcJMJOl+jXVaLlRSPZyoCbkZishBv0wJ
Ao0/sgqR25CsTkD0eXW35qEucoDVL9VNnTR8fYAZWLJ5imHzE+8kBLQDl1KfJxqi+FqpqTOfXA2t
OZmhcg5EclH05nimgTBD0cQdTfI5HUbiFmEMjtq+UD8ABpB34vJB7xiE3EP9zrLDEc5oYS7QMJEL
yIMTxG5wXrE5qDjo4WSbLpMdh8QAmWxeMXp/SqPMkeBG8r2XD/ef6GBtnJP6q6BrNaodAkCxWLK2
rCAC77fo/v+W/WQRC8YwMuuxKaS4jPQrnos0FEqh+caYKpKhar2fUMDkD7FH1hFfNnelVmlBQXza
m01ratcZn3A5Pee2w9kAtqdSiHXRJJz1aZPm/g/7cjCmgCd5B/yPdt0tiLYMpp3eLBqtlb56Ved7
vrfkXhrF2Mo7qDCXqI4X8T15xaMoZnIAJ3mLngfAWJolBQMtudoomGilvfoC/v2P63gEsJbLFRjB
Rb7jWa9WBFHqTS+TQ0VGDEk4LGEmGMjGD3HtDcuTqAtUMVED2nz9KNqDqxx1zTepfvgdzwVbtJVh
VbyP9nZpuw3o76Se0uYhv/dLtbJDps+k8dXnuyuQuV05VaKb2u/JIkSlQIWokIM0xPvvYc2DG7Pg
Kr8D5A/lA3/s9fwAIZIEGiR3hvPZMdvgZSJTKi3xs+CTz6jTuDSm3Gl6aFoJDNUoVEYUD1pH5lIS
7JeCQY/FqP2dKgPiNeYCXHudzL+gKro0kiSIfmBWDM49CU2bRbgp8ucNzqYXGKKgLDB0Esm4WRq1
TIft0amubaw73OTkZcDf/+LfCji+N4RMMoIC/nXSJUIYcEYGN5Tiaxnsfz4ApVhTW5jNTNDuDvX/
iD6uLmhs8CkU+5IwoJdPWByY6h1VxFyuW61jHfEyZA00mH9p00f+1A1nhaxkg0Mf31G6r8b6qs6x
XzmUPy8rrwizWF+T9t043UlsGx0ww/X+kfSFCPQgW2uk4WazXG/bii880VoC87sKtewua4ufmwNn
VTh7UlxutwJui1rF3Y/Hu9q6XG+OR1L53WWhYIIPO2wkheUZiARIMtdLPCrtST8AEABZfMxY2FeK
ODmKfPq0sJvzYWydl5tdkBnMQFc3tan5pUM+IaSrgOp/N9cE8//8vadkJJ/aoDy1Q70m2awRnMgJ
JhFIlNoM3NWo9IDizcenzKMATkCokTEhlqjSeM4QKSaQiA/a+PyTMancYpGxQoTvcXkfYsHIdDvq
gWe7SpGG47Ou9bcyP4HItG7K7QyxvqFYzGFBDxySykB3T5VKaZnD3MY1xJ7YxpyjlyHu35uWz5mp
+QWuk9wxD6+mHDEdHo3qqvXiZt7TvYAE4r7pBt/Im21V6obhtsR2j+CthmfPuJj7TofZtMiGM/9V
Iyv7UUnXKQHlW8Nkkg8xo1u9sW6xR/QrqvP+8BJVa/DJIL3sG/bOFll7GIhCae3EtgMky9JHAfmB
4nwDN5do7JoPoPwPs1lp2hRukxp710obNA3fA5NVIyBaTAudmbCax321soVwEPkfGu15KZgKEzyR
ffl5cU38xjVAYYKVPEM2VvLaqglizWVwUb8/Bfi45i4TjZ/OqoNkKZxRsCHup9oFyMwOsGUHH0LD
fRFzjNgY7cq1S8mNs89yhypMW2ws7pgMPNjuTj9Su2TlIDptbghcstPlFYoRvB8A4/kADP5wqli6
iLVI4iy57Vwbu5tJZ1E28KlRFpWd7mZCMjkLL23mpYWS8TaDn5xgslaFuxSC+1lITe1hS+Zm+9eZ
q7VXuIKgKpsmzwUyt/IpRm/zZwawVVkGwF66ztUBidcclBTItYsMpooxHmSIRlqA3WL3+HjB5JVq
KYpaujqCQD5e8BiP+zwLFz3hv3AocuZPnk69VpSrtTGyIyLM/yl9Ky/j//IB0Cr5DqR7xnBpHiM9
LEkV46CYZQU9+ngr2aySjoHlCXWk1hGGgMtSzVRDAICblYVXtyaOU0IBEHnscFDPQFegJPr30MXS
cuTpq4RwhkIfHG6ym8o+ZIXzXyqLXnludBaq/0ChCGg+Ul45MtU8UKdyXaGknBbt15ySP2sVHATi
ABVjtyi9Y0iVVEUCPQvtNOgd9L/bLm7v8OhfA9qUe7wK5HNw0xS4aRRmfouiOxoL3B13IZCwXK87
JJKzG0X8QN1LTSjy65AaarsADD34jhpj2CGEK1vpves6o4Ce+NuKE2iKH8sUFzdV5T2k+YzhhFXi
q/LumkdanLWsjY489YhL7I54kS8R7jLv8DtZjCnAidA8nTvQZgaW6caUVsz0KThB28yjSYvdOG+L
IIADsJwLbwuuagbXhRkdntT3Pa5LALLLN1wLV9ysktHIM307FHHGDHCONUfDNJDNq51+QzD4Tg1P
T330+0R9e+N/OM5K24fmBuQWfJAgxqgQ8TLb3qc3B9js8pkeuFY9O65Tv6ODnkkQs31N4ZHHKs7s
95sdMt43WmuGREzUlOeKZnWSJWLAJPrfo1494UFLMz6vRZdTz7eSiidnefk3HcFWdtm9/u0wDPiy
68t93UmvtT/6SGB/iQ+TqkVrZ4oBwCW9Q0FboUhPab7+qpE2a8TWMdRDhZ9829TcIozCpvD9BuNM
R1Ph30qix+ngitWbFnT/f122X6U+D4m3Et/qkq0exJuodmRyGt9MthgmntZvilH0fQMEzuFQ9l9e
dIXh01rLw0czPoqC3h1DTY4/yqh0LK+0QCr181eqcAMiqYgNF0uURbpZ11ODLUL1bN8Qu0ikXHLR
nwbnQGGM/f2/q+SKeT2GpOM7R7nmxSfEjv64qFsiujIt3s+Od3o63l0ZAiWzS5otYb2Zd66jMRPR
NkleY9oByRFC/p/SSUTpzSLErFlaL/F0L5Yo7VWg8NybfPlSi7sP1E3z78qFWI2IyYbz2PPFkAgb
6F1B44wczb5aLrbLOFY6T6F5fjb0P9Tb4w0jWKPLgki0otfTgI7TWh2zY0c3HUt5QM/GVWcEY+mX
f7wLz/p5yDPIDP15kb+AjUZlKIRJA/4qw3EHVR582q21WSG0+suGXjufMmzdIutiMhJNLYQwhfHD
6sGLd1Dt99PnELOckqA/0bnoJeL4exvDuzrWtCoqWemQI1Kx3z80fJ8/9BSctbeEFaI4uuqizvl8
kQpFTdnpML4VECmjRFH/AN9vOxe7oRy3xHQKtbfTQAo8W2c//S9i0v94gTPRxSl80KF3nP2Imso1
wQGWW7C3i2eQVCFVpkYg4ROH3+9P5bSr8knKlfb6eiUCh94q5ImRCYkEpv7SpUyLcwJE9OTeRQKB
0LXg/Osr9cLaHIp09xsfMxl1lHHSfOwYHckmbE4MUT2gK90jppHYHX8y9A+7gLkw+8ZjSPYy+bQ0
ONQzg4jL1t5TC+A/lHv7Z8MlvTY7+szCh+I9ymmAzDJqOp45nRivtPFpSZJzxLTJqqxRz35mR1wJ
Hr/Up4sUwojYQj9QOHs93khYAHxRXcGK5pPxkZf5EJd1gOx4k89n8v8HJhlEO9ELzHUYsbVgfIjx
xHePnINWiH8ShailV2kpexDe+WuPulRARoyAu6yw/GyjyEJ1Gz4Qk9rjadr+GVzVr9Cfj1g40hoW
A3HwEbNl6vMBBubZoiLenaIUT07LgwqvJerr0uEapIohNnJnz9p87kkYTYK95r/Phx9MndYbR/L2
A/7n/EMZZD0SSC6vGOmPROoiG/zYQuX45f/lHt87Tg1cl3MRNrNlOJk53HyPfmV8Nne2vYJx5Xw5
uWloTmiPAbiGt4ErDuR9b9tymsapvPsZy9SfBwq1x20j0X8WYyRPMw9jUtl1yYa+ooYk1eg6mT5m
OLqPZAGFGFV9tdQIJFg8l2Jug8xUm8eIexfWvfGPkIhjmO8HlzyB4QGFLsMGWhLzfGJIXeWMY4t5
MdYief943HYNZkdgK/9vsWfUE/iGIvkjWBH1H0oqSn03g+hQq0Fvpl5qSbBY91+jEq2uIFasjxMs
XD2CIS1wAKRor0Ezrq+5PpQDxI7lDhA2gQ3ZeEAORIe/KeIXLyB/ZiMODP5QwyYaVBBzTUkJ71V/
QQgsmWAuQw9oDqwtYiiZkm4315hiyUCQRolcdNnISTwOrrc+Dgv1h+OJWkzX9bn8SqZgsFdZqAkK
QltJZcik+dSQzjEUUNA2nKJMY6tNc4B0AeoIyn7ExRBQSdzhz1SbzKNGTP1L4qH1z0NLXNS+nYok
oGrwtuWBx+0YjhTeR4W7Fud/S5RlB/tC67LMeRthiiNU+DKnmBQvKSj3UQg82qZWQaxnnPL/3lhc
pCT+l5RwVVuiIgy9nf5LK6zov8hskjiWO/Vhva6Cu6BghpLltL1amB5pnl5XGvs8+xJg+d6zEGSm
72DdhkK39/oXBpXrfRMlo2mRwBhDOnrkisXWiXMfOcGT1UOd1fYFKDYUM1pz9tiKJqXlsyeKIeDy
3cGx528iZDuuJOQArvMsP3dbbxEpb9xyKayTqshqPJPvd2HL8msgkDazFneCHenN44qOO31kAUmF
SXDLJfMzpjUn7SWqWVHcsgAr9bZA+K7IiRV3e8J5qz/KWorNavgasxIjnfq1F2isGELOiwCUHTbJ
EIQZX8Ccai3Qg5JMA3FkRRqAwbNuOqMeeI1rumXXdSNeIaq7lUqdsA/oKp6GsiIo/xe534E1veRn
lxmzE0s4U5q2PCDJ/0VUdBjqR9kbGFUgfyT7qW7MC4LuC3rndDBFbODm7tdtQb+NCtRdlMzkDF5u
NJqAr8QRKtGEPAS/y3N0/OJCuFoEEwhiA4OcWQ4ERO2LjKFu8pCq2MWDhjZAmzolfxWt5oCv8yST
QqIe9U4ILlDVIj6mtR9TJOUqwjmJebf7qZZXap6FNFLqXtp8sz8U+wrIqJpa/jyd2z7gmaCnNYR7
1BjbtGWtVf6LM7c+bDssZCmD6q9mtooNgseK9QARhCs3HwQ2WfF2s5+hAc/1xk+kJ7O2Nk4zBUfz
Cdxksg4MGpv0P4trBf25Ed4nghgCZbl6U6go+cPyHPuW6B626SqsOELVitqU6xL8lV9Y0HilVczr
s3I/XYJjLqQsJRPzjSOSa8jvuKpC4uATPZvWPr7S4Zz4UFwb88PsmsMNB65fgzHqPQuN6OA87nXV
pg4ibygxQ6MuZ5GkaQ5VExeS0bJuBTLexuU+o2oHjGMCdMldX6LLi6QEZ1HJihBxzPJp1MYYd3ro
TqM3fPkPpZAPsjS86hUt+/ApN7qJ2fXTPzp8rlxLI2rFZBI8B0vldMdgBkFk43qr4WdlbN3H6cTF
NHgqj/NqTxN2wUDW42EI6bkFo1PaqKWb/USFpXjlaOqyLhTiQCUgwNrOjtLagAtHIlbPjxJVLlv2
Pp4d4cYedLYhGPXfew9GC/zBDH++HsLObaynEsklBCWA5j9s8UuMdCRnjD6fsL2PPATEB/MW7JxW
05k8PLLj4TKVP+KjT4Tv5ocrLx9YMojeZ7ZtkTge2XsI2YvW544mq/umVRl/s3JfKyM1U5nbVzpd
BCsUBLehymOBcoc4YblQ40APPbWaGBXt+bv9jiPi5n4JlYvI3Thf/qAo2axKYa1DZRN3CRQYrkRv
QN/nVftcHKMzWJfAjUdLIE4EtiwkuMWhLobFTrub8nRVi2Iw7aVD242pmbLWS7PVLjZOEnvoiZT2
ge9Lv5YY9RnV1I8bQVmcyed851W7bUzxBMsWNnfk6pvGftvqqF2W1jjD1ZJrSEU58rzXzux3j7YF
jrAT6+8K2r3maEx3s2yihsyHQuDH68cMNWGRbxaf8eU3RRh0/uKmRMkSSH+Mih8H5Dbu9Jmim99O
FH41UGtmiLF9si6ry/stjbZP3LqUf1ttajn+5192CHCtH1fPWTXXfr0DFA5FI3mVv9h16TCqK8lr
6alf7MSzAhYo7uvqDLVFQax4FH6vpjexrY7DopNdGi5eh5WQgpmyeqZ82hy/dSD/V+ntaANWLzMc
L/nldBiP2W/FAyz2bkBYxJmYQxETuWYjGdu93aOXa9+Jj1tGK7TXVN534OEaF5LuC5b0MXeXYfx1
QvDTpEWm9A2SWEbdMZ2vgaI4XNqBt7throUHtNlSJbNxnQE/ZEr5iAf12AaKyicmGbRORw7FnarA
CBFoBDHGOCJhLVR/+Xi+anowB6JZT4nQulbLJ9tEjR+eUvWh/XWkAuiSFdYapzjwc+JGsCjb25iO
CMCroIUl4nXGKA0sYWFhwtNE1IAlIyiocHxtePXZTyTcm7n5zi15THe1hQSdrm6CMYesSEaWUuyz
86dnxvMHHqUZF2KqUACQfBiV5sZ79vNmuFjiZd88P+CXKdfoFfd2wp0ffXEo8ivsdniflbaoSNzg
2nTRWjrjyjA4BEJ/GtbwE8aBQDP8F81Wxmly1PSIQ2O6GkSxpBLbzeC5NKbBVM0fP+OtJJjUWU2h
wtTBAjo+05Vc7SaCKjU5kdcmT84+D+SX4jND4cuCQgvSfj4yXS8CE7hG97CMyT1LAMjTEnxCOb2e
+3J6acij+pg9rqM3oNpm2VLLsX0gUzsESsM9i3kPNPjXzmHHJdnuyT99sPWH41jqqyFn93R7xNw5
CTN3oeYC9ZE5+kNB0kAZ3622trKHreALBAyxBlmRLkQayssU2oP7dF9iWV7QavqAj1p0/3MmA5NP
SNWwPqjA3/gAooveNGFlRchTruNdUd3dCbC9Vg3UYcRmdED6QHjd3sXaGeopRqQ4dI2lbYYc+V6H
kTqFn/tvQSfEHRx373PQmphvUMy9aoYHpJ2+0/sUczdE9Yi+Es+rY2wvxszFij8OXf2Zu3kMbows
rG6u268PC7dAG+M101uLhBLUy35Wl0qTQnwXLGSo8axA9OOv+rWIG1nnNM50f5Pc/ji0RYK2Zlhz
/uUFRfeXPVtmE+Vtke2+kzRs11ea/Njwkn7WajNEDCTGOo7kkoKuO+hY1X5QE3pkrNvUV7Gs/id3
AYNGn/6nkkENr4hOJ88Q3SsajboXvIG/e31yqd4+dJZ+gyayxnyvBncD4nTwnaNMY8JE+fnYiRne
GUj4ncywMF3L4a9+sfHJKIN/kCN8dewOUAYtJkp+ZyiZw3oMGOt85K8KzAU8PbddsrgKH/d1AV3u
oorKMWAQgTf91yGpJ33r5gfpv4pDzxpTykEORpev4LrzVOGRclHsTx9Pm0i9m1TyvOqroOH6o2ez
UggiEoZHT7cf1nzZz28rdgIKoGpYyJLVgtwla6vUoBwJ3A8IN3tup9s/WayqBBZfqmSTSN/AbIFx
zV0QPZ6dBB1ZgIK3/tHjNAKy21GqgoM3ZQzqA1xH9CcIUs4o1hoGABvtzo1esbdIlM7L1cCZl1uS
DlzA0eE8xZARw3sVFmoP82NptaEn/IbjlBhuE8C4OyRhslqGXt5c/PAsl3LvFQdu+ZHn4G6ghEkt
5/6/eXgsbHvus5mEmkOQsBRPeqbbq3dqs2KUyKmLwFP0ALmA23oDaW0JZOC/ApeO/XH4jTWOCaF6
kPA3PnIY50HnjqLmQwnRM2CsdVH/54nNiEqhtulSN5ih6wJEC7ZenQr4A/hvd7Oz6UjHBnnCG+mB
asWsKdw0pKud0o94QLk0Yz6HOn8uu/rxsWA08i8p4NnAdZdUOMVePTI2+WEOo6BSjlK8SS4b78PK
iZQ/FrzLqci+tJMHDTO7GSa6w5S+jtbPKjCpQgTYs1nt6IQCAFkJGYbvCwKHhOeWH3sRr3dxLgR6
gItNyIQMvSvVSILBnPxuj1CziTBMAXf5C2swnuwIFOIhOQQX0XAapUR5gs5fqAVF76lMdNN5g5DY
GDNL57zXYJtkYstkbVLPyIrdIR+nrLO0TaefL1sSy9YRyqemrMHxSD0IFIak2BXrDTLxMVKfmFpg
rQUlnFE+J4ATEhJ0WB+dqJf3+2BaXiOuJWiHyr9CqkLShQEAzO5F6cYhE1UyFf7rHcyDD3FPB+ln
0HVWEVqXzXmHmg8sLoT2nTDLJQNZHSWbfKimopK+SjgvfOd5voncoSUvu/2IzdlDbRTyEuhrtE3N
f5OB/LeKxmIzNKFYJ1BxRA26Anvy7/+BRaZJD5tGf6jGGHMigFVgGuwqDTgOG/2k5g4/Kcg2QyGe
frLjwZUuXsQEHlVhKYeltXVLCzgY+9J4IclDpuxAm9kYsFO5DZALBhgUcb6Ru754Vup+Jl1yuzXL
5k+2Z+64d9BzzBEvIggpBLpxanYhqJZ2yS4aNGCZHnA7EK5knbFcFcrGrJYokTcvYFZ98J338ucm
usAN4o50eCfhuYMl85FZqBc7Da6Qo+aWiS+wJUj1qwLIRqoP4nBlvj3TRO81g2+xJmq7BBEPn0gI
wioVcCvV5PLnUiujJO38yy+DCRQtyYeAbZmzLsdgtRYaaHNljUi+5WaSgPQUW9sQWKAKkF9AAPUw
uE9sEhZZ1LqO0sSjKZiNz+AxSrVQW8vqnzyEn22hGCjb6M5cB2tTKw1dutwoShtg6By23aXu1EHd
vHbYil+DX7BZLAs4Nb0a9Og9LUglHVVwDQVQxZbXhBlBLH06U8RfcYuLpB5tqDVjsG8z07jX3QZp
2HxaRECdk5Ans4j6SqBE56JliLTn4sBYHJb517HUPYAq+nCiwYxgwsUDnXHnYUYzn3Y54OeQz+3F
UbWinr2r6+7wpCsFaVbc8pNJus9lZvgMkKwx57y5m32At3Wjgd1cFbfbJGzdJzUdzpCRuBEDunj8
g5Loj9xWw9R6zOgGPv1e+5EpbOnFIk+89m4Ki67cNO1BNjI9QR1oBsJ3ix0yEVHcoyF+KIcuWloL
YsUC21ywbDfB32UjjUTgesIpiw6EQjsx4qHq4kDn8ppYk+mccrS7/VSQz1ZYopDyYW80+BmVeOMS
6m36dJvxf5v9jugvLbPORQdUeA/f38aNgqfm+lp4RNXu/CtM/spsXKJNcM9tIXFWslSBXhGYATaH
MxWpO9deDXfYyUneGS/96gBm891WAuukhZPHUH9/5jsoulKyCziYfmNDpbA3xZIzZSPIrudbTB9V
5u+BG+hY6K/XS4SpKpIv8fm1GGnP5Gq72qr6QjcxENAv8bsAjGIgV7NRay5KXS5KrxXB0NoASQBf
QFVYbK2NgPcm2ldr6tTOCdDdldzWIwUaWmErqbJM1RVjUn1ezMhn4VSNY5HyZAB/Ks6hSNpeX/JY
8yrDFUji54j85BfpRSGUHeoiEHn41wsY+va6VwHAtcsdULhqWyR0iQAieWdy6L4XWwhN6h8bDGqS
lVjcXvwk4K60iYVgxm4gpBbBMQXWjKqDKgqIbk+S4P1LbzpfgeL9YtYyeALdeLyIzjKjItX9hA06
lOIPoOHbhEDunE6XMhWdDVK030b71U9AIzgz3uHcNgFdQCNCPNljlaFp7OjBO1Dl/H4RUO3PbI/U
+Rdvc3b6ijocv1nzoW6ECBNqp7vJux6Jd1Bc/ylXkz3JqFKqEqy6kb5iOdxHD4p7m3MJD0GmHRti
8bAgt6gt/g7ddiVXwjcYrBl9l2Fn5BNWVjvhzkMH9Qj3RO5a1VYmbwFo1+JKKeYcAf8+UxsxOOEY
zSYGNv+Q7b0nl5sSXZbSP/n+9D/if5mata6MWE3wYb4g9kGcU5c3x0VhBU3rxgGphWCpfS6JQcBc
3I087LdtI6sw+1RiAfJP78GY3gkjHK5t8TEcFsbZ66Wxlp0Dgbrg3w6wUwk7sI5PPZ8I/EhpB3KV
dOiSi+KTSn1zOfEKK7Xg5V17h/vo93iLroKjUV7djjO6XIRNWneT1uVv5LVii7Dbgtz0UbmB2tum
rMb/hNVaX4Ve+Isxs3+RvS+rdST1WmbJ3k+qmA4/erB0AoHeeBpvmIygqAC8ZDKj8XHHuSINaEvi
9/T9uGKqH4JykdgNdFhSTOU3RntWZvwi2la0ruubzbJHIulgtriUxwrssFU2rr1xpF1K9K+o6B4a
V0j5bhg8Lc6ExYOBl2u7F4al3FlTd3A091yMeJFRQiWW5+T1PRlrbOv6JWcxHDZ4DSlWcwuL4eg3
rZqyyFNlm5qSgIeC3HgFyBOXRJWnmN99TCxxfivNmQ64Bc4VjzDI4ppr9xdgjGeIClVItTzooacZ
65/367NLKdp4jdQQweiTuFDNay+qpPKFDX0Ks9ygZsJcn7YCu1wgcqa4dulLoEZ2Fo12HHTFr3tl
Ds9+VzKkO+1h16kTTQMk/ziS+n7nWNjFBVqDuFiRKnvBPEsR6OB5VXUYNFM2wCxAdeXp7qEob7UM
LmTjWCMSWLkV8nepH4Ej4PKhw/Y5//JYGVteyLsy3XiBLwjxKya1tSS+jWEobehdRSFc3poLnE57
3fwLQGUHdUeZ7/pGkymiD4X3+Sn/ogTNm2zMXHJsKSthS06BpUsKBIWCstsPrf33sTeL/gtEIGdk
1YibD1tOXlIwVBr0DT+anTC64AkCJP2elS+d8swKoBO0oxAmQRAe1GBl3BfOPoTgJRGwxDVOWLku
gacZTyzvoxLLCokp3iytbnv/adHB7KaHcUuKTL97PTAPkPc26FSkXP1sPgRJ3fWojfI3/0+Azu6f
PxoAD0A2dejeg1jqwtFIFVI3aSAN4A7p2v9dI5mJN5KmfrWdCoocNmpDKOTNMQwJ1QxifT56LGSg
4+ViKMy8EZKM8uzteDDBdMVXC3modzX4YUGVu7MocjSYpn2XSwgRaNvOZzbgSUCqBnW76XweL4Xp
RP9VyQzq7HjpEt2TJKdsmEuHOUVwg2rUBzIJ1iVeruMoK/loUpjXQ4fkF9XFGno1zKb5CdJ3HpAT
IuCNRWER1sAOhYXsji7DiF+3KTsngzVcfMl6SwdXtIyKO51rIwXk77g/f977vVnKemw2hge/Lciq
x8JWmyjoaUzNnTUCaHoURfDbC1Wj8q2HSIrGZh3RVR3LwtiyuyC316LG2x7EglbW6LxBIGAPzhVz
dDdS5Ch//DibO18J4d+6zvIVw2Su7otq0ogXGSDDTME7wmzTs4htxYl13rZEEIZlCSDCKqJRDBp/
3CHsMU4o/W1QU9wayvCsu8wmtWNyU2hBz2UIdRKctzvC9vB3S69PfSIqOXLthAZsjdQ811XxLVpN
b76cnncjZf4WEWI8epBgEonFwt2kwT4BXBB8PYlavo2j/KM5jqQWyDwayPaOI1VDq1Gm9ZqtzXNf
/ow05FOlba+8w313hSQZHyaz8dP+7jqB+dCzuDK8z6I3Swh4nbtzr5R9ZwyfjydPEhzfiWmt7Fo8
K+Mzn+5k+CAMD3qyvKtnCrRbvvQ8d7NKtdcUFrokINFaFwNcT7pmtY6u8a4Lz/oXOoWsQTnRKGzD
CFOBbLpSfoi5uFv+5PAvhphxHJF/TgADSRVgyLYpUxZ3U8NQsVIMdg0Tys0R8QkWWOZ1h2xc4zar
REOjI9tNroyJy9XyIscViRwrbAO5aYYV8y9l9wGeEnRXi99al0KipWJFHS/QWxCbW95EW7r/G8TF
ynZiHDI0gZT7B5FTTY9X7W7TuY+ro0NyXYYgvxvaxD9hyWZ/GvPzfzkjGPBFDBUOW6udFj1SSZ5u
jWYSMrRfaRSS2gFUORIT3CbS6W5X8n79+jM+KHoOi/tRT3iSrksKBL3Hai/8km9r20n7B//+7AJ/
NFTarjndbR98eGK2teb3oLocg30FxyJ5BuA+c8GAvERucL8XXW1As7/OBDIK6mN4bFS0q1IY2afp
TusKSCJTXB79wRSczo5Pc8n9V5Iet30/fX1G6GDeK8FzFH03xliaYtQ+P6aEaX4s2meZxRkZUzbn
IXP/kOHTyhcBOHL5Wd9dldXg4L6mLz62kNbBYiaxqMeViHwwE6i8kCDhz6P3f+/+K8LhM/yLGJQj
6M/183Y4svdEzh52mljSy1U41izigfeTXT7aPPdHU4DZ01ON2GGZNrEri7fLlijaoktarVP9chGk
Bbf48vRIaLzSHV+XYoiy+2PDNGnC9XU9M7caQI6u2CdfzP2wcd/m+wbg1J/d4HcaIo2q2/gAGFYM
hHwMRF4OSdIsk6Mj10lICte1uf3KjQJhFLVUSZkFmO63kpEizMYbNyrym5RUcqIUa9rRkjGFShYW
79y+kKwEMYVwDYYI6rc42cmWsojEJgxLyUG7PocYO6lZyDby3FbhS30X1cG5LvSnWAIUIQs3+R5A
Elmo7x7evA4aSGkHQB//rC5vDqd+BDh0yL3TtZcupn+hw4H2nfUH+IfhzbnnOPwUa8KDliinVv9p
bU+27CyQAPP0rYaorsQBddM7pXNJM6iBvw//3SBgPaYDsr6wpjDraipFXYg+9hRnT5pE3xmdrQx0
piskaXmHcC4Cw4OgBF8MIsYoblO0JvNGAAX8/JiLUG1unDcvkTryo+2aC6EgjIiFUcgy+DIMpHXj
uGH/2hDHN3sYtVVasExZI2ZCRALJ94j93xv2IfhV1KiFFaouuIL8XR66nK2bBCg2NHLLlLnKVqsI
qxs3xSun3VFLh4yWcc9YVfLifl9WvEB2sq168VSr9H+awXQ1rINGU9q2RFEt/MO7cJKOx7QXGZcK
SrjJfi2QG7OcWfJSFJssmvzTRj+JyPmdpooIc+6aWUgbNTJL90rKNGInR60Y9uh36jyAcFvcbobv
8CjjgSpDGRL1DbuMecXwv7NV+Cq3nyyXY2/CmS3CWfXOHlgj3+JG2Gt/+h+/0ofQ0g75WxHkJUZP
kp051kotzXvoWVSbO8YQQCXxizPv/v5RmsK9FcYyLoAv50zNW+mGY123zftyDS9BmH4hgJMa2r7X
ktjnU5XImVPVCIQtckwAPBspkl0U1K1q5ZUsVdwgruO129GQ7Zw7KC0KPh1SwkLnChiP4F6kIEfk
QgJmWMan/IbmoPU17BeWGwPE4qSemgF5FILzcH9hd5vfIqhvxm4YvBDyKe/7/E/WuxW06So27TzB
ULhQw+XThTDkXADY55uk9faji+X48iBr6vgA6lPa8tbCoupizsg3efxzhz4RTypuHSBiSoMlZkF+
K6L0or63OjyT6y5MzEIzZCT3Eju+sV/6Bsgtm7ITnZ5BQjC6x7sfuw7DAyjj7Xla4RPLWwv+tWFU
/58RvYRCEFNkUNqRxovYAxtwamtf3i/NnBr+ooNIfvxEijL/kQQLYL5n/2x5BnkzJ/LxoG6KPYTU
QzcbBxOgHiTxQx6Njp6O2ymb2Km3XzpOIGz3if4MV6M41WYqgOogtSS2wDw3J9qFBmW3bzMCCNIK
XXUHUtc3UaJJKWrcsbzhiB1yoaC0akVy6gZLahSYgzSwDWpCqwI++9pDSYd/dRN78dFRe6HexpGv
rjUtWi5ikxIVgrrjFDuD8OB+s8SE2tr3G6vxEgbRxVJKDDofzdC9Ik4vqPlCQZxFu7G4kwd06SE0
wE98q+TXqt2eIhQfr56iVpKjoNpFN+ytoI54ZOgjWJDtKLbV6Hb13OVmx7iDsbbI5oktomtjQ3Nr
9J6KTIAabpBzbky35HJqP/T++1DLeKiThd/tTq3uAHFV1etDcuaeEAMtH/YQIpCMLh8ydnjQ+WLA
o00zZyl7AQtAeCKsIhhtIey+0BLr0nXxCqkwRXF2S6vQILQ1hh5PD5VxwpWfboq67KNjW1jFeT7a
EVA4GS5hWkyDRAChP0B3Q09XgB6z3ey6F5RPO0Gdk9KzXGLzv35VMfaNeFbZFO41oy7FIFodxqzO
5yFsaSzJ98pSUHKdI/MeocA8lzW/Yt6qMSQfnro02NEc0cHGXaTIesHFYRW9XN4rb+tjY/i7VjrD
jBTiIZKODwZlAAkOtPP9/h7g3XKgTQb4KEIYeh43FJMM2Bpswb4PFQGF1xww1WVAHIdaPmz+2A/r
mRlLFTbSKpRmJU9Fivw8NubVau0HevyElRHX7K9vUBIxyL2HAxSc85bfOJ1htw6cTluluOqEmhf/
XQtBRjJAG62HUIcjV2w55n8voyCYBKC3s05BiPbUQsS2/NEsXVWNVOVlAwZUY+YiOBqZIIzcwJQc
l75N0p2hk0KsfhOhAyLp668PQ6UfXHskpT9NmkrNT0BAEnWqmQ8SrDDVTo2GqZzDfGMSuStNs4Z6
M94Q3/xYBCuRdB4aIWJTXEPRo4NXk/j/xKd820Dp+wtQwkT8DaSmj3MPHjxj5If4FDGs/pV03WrX
g4Lr3tyUjYgSjae+pDNEyqyztHdZ6h2OSKT+n3bizTcjkRvMXCsbdMvIUpNUwJK06uM9KVTqIMmG
FbeRpD+1TD04+kWQHQymo3y4thBooiav+O6t96UPDpmvE3YM4ddD0sOrPlUTxqqb3wCOkmgpMzti
fjJpIFbS+F9CUEmh34OpxWy30Ske/RdYOx7dDtd7sdn/cFiTJ291/nP1nymrAzbn9xnKbf+z0JuF
KIhzdG9dtis2O72WsXjLjgDL7URFO5Zc4RAS9lwQcUJ2Oiez8+MrV7sLtIZVOeRt65Z35x6sbg2Y
YM/2mqurnLihwYUFKPCm4vsB3rn8UQPph6YL60MAK4LD9N1mFj3jPZqb/fsPYuxt+2cpPSvc2Dxl
LU+SQP/EJmlTOvwKxqVFNQUY1pQMaabLhTjbhYydJcy4R76has7JoZXIITZTh7hMjLwOHWWfRKWK
kXk6gSdql483/CUvuFuWJDm+XiqcmQDlGVViRmqLCP+SOT3X5kbsyZpHvgLxKBdB4pnygH2TXTeq
eFmmygRt/bH5nJaGm7qpwnjIAgu3rNgPrCmEXs1A2ixxtG8oXrp3MFuBh+yP7TF4KVlQw0hHcL1q
56CvMftil5i6uvS+pzjBgCAW8hrckD+QlnuHgp0yexkYU5fqavwVxgoc+Yk47SMynp5PtUBNBjsw
2CgwyE8lJywaAfxQVICuNUoJMiWEyhTQhggXymbM7FMp9G7GUt5Tcv0OdaoHSgsLXJJ0NHxlmUAX
LemSCK0ywje7NmX3E7ceGpt757IUIbHOMrOvR5IQfmQCNL616kdInyvjLxf+CTA6PGVEiDRv/4rI
iJ7l8MZs+dxdlshdE7034ngcaR1z4NFsqPH6Yvk+3/BMMvaEEV8LP0bmD5mT4krTTqEwdkFZQYmE
lK7N4x4u09yw2zck5suhch98gfN5pCRQl4/NPBpxesxAF3OrcUeT9rRQ+4Yrg9XCU0S6rVXiuLKb
r21qy6J99mQI2poUmFc+deWisagNP4fKsZWmvGENExguymjFRfAUEShmdDQy2r3/310qPUWse7rz
VdD6AD8YO2ZRlDJZ3xVcbHd32iiZ9sK1SVrHT66GrPpaXgH0icp5j7z36aXh0tJKbckK5MJga6tJ
crB/vxzw2JaQ3daAzuBJWumsRfoNIBB9W9lzYCyclDWOQeFS6aZ9SFdbd3FQz7Zf/ilXc8RPgQg+
PprOFvhqsduUC6hrEUGWKABfMHrp5qnwUo8xscn1tlduSOkKud/12Scyfcehymx/xtYLctFLsZkN
kW1fQDvsuZpLacFNECbQdu/WQw9pxKPv6J32asvanCPzjoPU8ZcO2qL2cm8hgBsRemD/941k8rAD
X8NZZ3PkZrrS+OTzvIfHNtCdj7Dxi4Jc++hDVOFMfs3lpd8uEQyLvBujvMTTGkS8d94DUNtadLAH
0qc0dubZ/eMbu38kZr5LLii7NYlc7g3i/EgEvG9TC2wshKXTg/x8hUgRFYrevYmz9F99j8xZMp55
8DZBsqA2u8Tb/5jCPg7gkdUfhaZH5R4r1cOdu9oHfj+0o6Q1Sm473xk3gFzfAwIu8hqFKMt/H6CD
jdt8FxvGuT2mzyEdkrVHrN7PJxPSj/oYhFijziUD47kMZXiSgDqXod6SrO3WPkTu34uc+tiJZbK9
3uhebAdIpyuXEh3p6jXA9Y9wvp7Q9wubwje3U+TFyTebXfFavnur7QzQYG5Z8QEkDHSXQtFkrd7m
oSVVsu1z++nKNKGMVPyajWvyLKJp4C1kg+sahxXxZqpoM0DzmB/cLAOrZw924dbn829Gx8sLmhKh
eD/t9kdYFQW1O2GDf61nYTdNqiqB3vSxzgWevIaDa+E30lPH9k8wWTPxEUGSBmf1fyJSnaKbDEF4
I/oeeNHEMCr+EmDmwM1NJrAfP7ipE/vSE0dA+HII9nRBkK2Q7jJlVzPbydflrT3hzCfx5EVdj6FM
+eYDqmasCiGUBtwh3pcpoaU8jouYzivJ2s7nVYySraeGCpPpxKPxBy157UWLwhIBqCOpWuKTYEks
lsM3NSPa3TUscoXyXWlP80GyqOqoByWjUOoZ0+Eb0tl8CtadNdqFg55EaOPBk49UbRNtyN6NaTcQ
J+2tlbo+rSiXHRhmnuOGgpaqcXxA0K8Keb3sLaEjA7aQpymoarDBE/X0xoMQQ7nkeb+l0dV5pn0X
B+qz7HjJhm5f1DzFzgcusUxL0h6Ke/0Y1Ihox3YLytShj9WLcb/EIoAlC4jMHwtOdXOd0nTBJwx6
6NOACiq4OZ2j78SX10kPBuoetBLmRboiswH1H8D8TZCLszac2IR2whuzvJvQ+0h+wHBXkGEMJAu9
hXnTIKCY+m1jZvl0zaM+yMFM5z9N6Pr7VeMM3W8/K3x61pJekyq1Sz08LIDdRagGh3EaP5mHkS/b
b4/Ntt7TfpUNzW7NN2aHLpCR12OZOMN7qeQb3a2vP2D0gU+q7MBN64n3WASbEncLfHDahScsJIkP
EYDKj2PHZpgdkGDVmkimCSpEzEUr8eArpGQ/kpf/TwWtgOWYCUZLRtP1DEDumKF4R3LU3F7XcPbP
MJY2QZi45egr+xSMWVGoyWw+Bk7Kr2K2OOay0YVZbcxIG8pZ7FiXafsGWuC5sITFKz1v1JNeJ7We
bfiXR76tOunznuBWGNLwi5TYShu6RGANQqMQ2XLHlpG6SrTA4jNQ4JN4nx2fs7Khdc3zXW74wo7Y
htLwKJzbuGPJrdFSwiAfDDtg7BWQN2GINpvMeP/ZB/ZLxQs3pESVq0WSf3BJDAESn3P3L1AyXgkL
CecwD4EQk21Sv+nqWiu67ctQRJmJictcffArrd2S0GEHVJfxv2/RTRoOJNsr9of7+f1Aqn4Z+nc1
V+ZgyKfojMGw/AYW7Sm4lVReLHmy4ZOwSdHTY2DTI41Ua8llIwy5rQRYwzsIE43QhxUm6kZe2Fux
fQOg42u/SaPBTYRcTVLAh92lxIWUW9GS4mQkC3Q8cWNp2Mz5C5Jqwi8cF4Ko4eIyfuVmQm2MJiGm
D/Cs7eW417CIc7rQkFVGAtJn5+PyNuO5VVtmVE5CLQoyhf6APyG7tc2a6HuNISu4n64MqtbM9rSa
z67TB2iT/JkeBZPVZjUsulZ49sSjjtqkenkm84isYP09pKw0wkPy6Uxfm3+hnahdvZZUP0Ln3z/2
XdFL1Yu75Jk9GlaWymS7Diz++CqLFE8BuyuKqZ9n+BTadp8nBXvJv6p2f2lxsW8SfOKz6pBam0Oc
tmSQZowtRckJT3y3tzen4n3r6XLVva18/CVGBTBnLrSLHRLf0lFoGyPFne7jEV0aiVEm+MA8sF6Z
9mlzKiQq7G5lrsaeM7Oi5uFJI0FTcGVmoenZTD2Fh+HIQJXLJGLcj9E271CWNpiZ7dYK/mY1ZDDJ
NvbnQ0bYQHZybQWSnijNw+QL2yDs+fBr8k2XUBWPQhGR7NyWGPqR1o5ZAhCPg+T3LpoyIZ2VearC
HUiRs75TuJcteC76xc58ammWpg/o2ZGVM8FL86h0/sYInftxpG5mSrmOF3d8vdGpnhUuE96e68wp
JtEXKUEWJIRdgjj8vL1WGHBulRaRxFPplz2Ocy9AL2/NxXB1xOUy6eyVR5vLNz3TVsLE7tQ9GUpI
96h4hB2Pq/OaT5J3hvz9UXJOpO1KIMMR45jUMVqW8K/FE1nPSai8IIo/XiuaKlq24JBsNWdLzrHh
3Dhh6QmPAkouUuG2uoa3tk+tJ8i5kx+NMtAYpL0gcu70BqMPmmM46x37cMzLtXUeqRDgjJCuQh5/
FT8WUjKKDJpJR5wptPwHdaagKs3nQswti7GpmiRNUY28XufV/6iayUOkCctXruORaPHPoNGN+cvZ
799VQJ9tYx0WxqvSSfSq6WcFVhvdKE24ce8ji62Io2t3SjqyUouID3fujR5t1zSe8Xj1z02ZZtLe
ZJCDPtf+zkvBRZwjnWhFaBGwVQ80VZIVkJqxlG5MQgxGqiDlPrcalMJNWSSV6kBpobdcKfVFaouL
rg3bGIx9291uN72aidT5bVsQgS66OUnAHAYgKqtM4RA+hqDYxIVt9IQBedEjph2Sk3Z8Kah66gz5
CYoUnQ/Bq873JnGMZ1qv4L8bHRSs+gpgZ2tEdi67+R+vVH5ZA60JEh5KyzA9+5FaTgZX5TsHXg3Z
7jqsE/3BTpxGTPBZPD4mAJJONpjbp60l2LN2aUmI/mppGJW8/7GgTGiH3nRV/IR4z91IaF3QXH4b
D6bHlBwb44PZ3u5QWgcsm/RW8DR8VqeBfowHMzakaMJ5oQj+W4+vW9at06zjbw1cCNwqEB2IN+ac
dAF+eB4zeuniP0tAHPR2wW/vYgCoTTYAUtHfaLzBjT/sS5TqyIfDq5ESTuITW8AtVvw5okdorVOm
DEC0JxGljrNEpZuEXUI8UYW3eTsy1UrG9QlzEmJLrIQZJEac8Sp4bb8gNMByqL6rFeCfkkq2nU+c
M8ijf2fIm1L6RNpc2g4IwSMvzGhbUHvZlNAt1pxt5VswKc0xguzQBPsP0P8XYx1DoFcWpCZdy93n
7ZeaA8A9u3/JIMcog3pFA+taHr2oQiR02Z+agsbRSHJazJS5gQKBRjP17P7bcGXGYLSMohIdTOUu
BERond2KSEthXrWxeA1kKgWJ/dpAam1Dj13g1Bld1d/a7UdgUpJVFX9LOw8oz68tpSEZzZqYuAVf
WszIRalCJ5pWEoICaNbhq/9TWJKYwVhijyYhiXN41a0SVJDuGIxE2nNTfzZThe/J/AY+slFlOzHe
+dkdfwfYD93ob+xMGFcSBHupig57H3RyEMr2mIFwkb866cwzHaJSJCt3mZRAVtLAD1UwZeHJTMEK
3feLIXg7rrjetqKqCD87tjGrr4B1wmVWcozPrTnZL0k0vk/dcITlIe3qZL9uzR/0infuWsPJZWdZ
ffWfxPvJHjanO9TZezijCr4Ur+o8STPdZvyGGulLUUJABnhG3IDJbDNbjXtSZhyP5wiOVkPnLyhM
4prwzrvYANgLyZ1EeViBiLSciG6e2KI1zOQweoo12KcWFvgXdYjFDFw9oXEFOhHXZUgrCMCaTRvY
LpmteUCkqPqmZB2srZm9MKdeE4V13TY37WCxJAlDJPvmZ5QifBgT1mDDf8e6o4ALG6zA3fYOm6b7
oYd4yKSi3xsx+olUksQOCe66iwW1K2s4E0ly44xagQ1Zp1W1erHETu+mr0m6Me/utrJjRMHIwHOS
2oebZXy63ACApMBxzvIrWjUYsqv79nllj+ynny2hJTbIox9GQthbWv0qg9uH9+T37u9hpud7pgWr
037cmC8Kazvw8oc3RZopEE3tuQ4kJKtzlIhhRVk7wb3rcf65o7Hb+keSpXwqb447+WgLpvBeQ+Xf
xFNCntzj/9KjlcEa7JGR+kTza2049JfJcwWNgVn32DSu50hhXZxrOh5IRGwsFTH8gMk0f0/C6ol2
dSlchJsPKOMjRI1XJcf+SbYxbq3ktJxXJVtl2R4TsDdYcpdqU4/8ZXy+TJIYoKUElVx3Yk+eryTI
yatdzt3roS1KglNF2FT9trfHZQy/tdvRxFjVff8kvzEqcmKNTFswWAe2yOe6VR8ftm5igIz45jWL
4ajinjFl/PN33kzn5WlDSmMHJMIJlAgcAlMcY73GRpnaPXuvg5LwlA0efHSX78wMp1KBDSu645aw
ADOLLsOeP7cROA5NMf5puF9JpbAEs3nxRi48inIVFCjxf1eHKDSJEdlaG0gI2fPqtFA/ytEBoVic
IBPl1yJZhDijteh1XY+OPMeXWypXPmhFyytLUBjT3UMeQKmdHgFLzSZL8a8yxt6QE3U2o9qG/bYc
8+fV4Hxjt3h2AAnwnQQ3Np0UFUA/VYjTcKZDBQzTZ3K5pwLGpJGkTKMHFrA9JbXr/oduMbNdrkVV
sB+FheLelGoBaG9Z/skMqzn2uuZNq7ITJbbgPpGEc7Hxy1uuigWrPlpEgt34cdPoNnPz2rRowgjk
I/zCWScctEmn1G1EGl3X6RcFtxDTZhdvFehRvAdY3C3tOLy4qsVd1bSSEnZARQZj3+yrPfm6A7A9
hvmAogPKzK68ngB8MCk3Mru3Qr2DRrCdvBcNpyXxwmE3VfioNesUFh/Rt7IXVnu5pE968XQgUtpi
8YNTyI9qfcpuvjfDJVgK5wucz0hPw8CNIRH1YZoJ1AfJ3M2c+eQA+AmNIIfOgtNnyMiG9VGITCNV
xfdVVI5DCz/JsDeB2fg1Ldirzya0mmcRkhrDhMcgkw2urmLV8ZEksV79BpAQPibHL3G4nCUQHQKh
0k83jcY55qEHwi98Mc2XoZ3CcQP2yf44gXomN6GynSQZm+i8Mj+ADTxaKi6FJrPnImSLZpBIZsaB
Uyfzx3FOK5HXSLjb3L5OcCCqsu1vjkdn/dysKOFRkdMcvxqV4PmN47TZzLEwXKQ4GPj3MabAIt1v
iRUa/fEaGJs46lTqWhTuuhJKfrytMknXSJYPxAJFE5qpC7YSIdpZJJmQOpxxNpxuFDN6SWqlYi8M
7+FX4alIPk7YQr78+RKbyAN7KlWOJZOobZ7EUwlIJJn/ShIQddL3ak3q+RbnmfBv9xtgQxSY0c6E
D7lz2EhiGsUFUY7U/gTiT4x1HkVdERgnA26AnVfQ0+qBu3DIa1He5z4QSo0DjybmpZrI5ivCpSkU
vuu7MesY0XKEW98RqWKyLwnnjCnpl4VDS25AgYzMaMx6mmZxlY+1UPmEDi1zXM7v6u9IxlwopXSn
gYM+Sk6FR87ZpKftpMi+9xkYeXpm5sWRRxCLHs3r7NgPn/DW4GAvp4u0R79rmu/du/65/rlzxzYj
1FCvkK+yxYnwWlpgJN4Dmpxk5jj+e9hP3j7dIHJWkYOG6dBx1NfC4Enfc+bPoRqiebYIAshzPUf7
sKn9iVu7Js+T7nfB33JqJIFLgif/WTzr2NVZxEdOXfvptzh7Xynj+iQKBBZVYwnvxJCHIs9dCTad
OgxMVv9zVCrid96l6pm9ZeOLJNbu3CdQrs9iU99Haz3/FJs8+Z41dDwVddjkqtO8oGbbnaigvtd7
/BMG6Coh83EiIA4QUgJRnZVFQMNHh5jCujl6RzFmHM7v3PKj7VVRX76WBT0OS9BW1vJ8a4JEh4mo
d95SA9D7DdF+WaCZNEVkFRm4kFovBxbV+/SgZLlNQ/pl8nnOEZ6KKX7Yp6UjBrdSS5XdC/YHRQvG
H+bQl9mn99g+9TP4166hZP2rZrVW5Nno1cAJcy+nGlYfBsrOy+QOaQsFH53TVbiY6UubAj3RZB/p
/JiM78kLwLkypHi6hKDdpTcUoVDAb4d6ggiw+RTIDXLhQsIV5viVa92MCqQWc7YM5s+K4RnHOwJk
1cglV23GbOYmN9meibqfEhlB33u20YAsmF6AaqgVvcvgDnAus5Kc8PvzKQptexxaz0FBjGFnLq++
cOHiyhZYTISVPMu/4aMJj0oTHucPVBT3PkUvOIWKbaTgRaEfTvsimFx72266RgoHz1Hn8IYzhn8U
DySfBXpSQgdN2q1J8dVEveQgPRMV33YnYLwUu8+mmqrAWTRTMw0MEY3DVwrTOBkU2hY7qQflXgdj
fcd8KqgnPDF9OU/LGM6creF3f4B92dpBmnJSD+sK6QUOz15E+agwjI/JASw1pEnCVmuFQ4XvvPgC
Qj4czsXwV97YaL3EYUh/BqtgDiqo5RaUPHidwSZdy8xutiFBTWQWfmT8yKedI8NN6/PeBlPARkpP
nZSp6kUn6gSeDSUs2AdfDULJbtsHImw2UvrzwwnMc+8Egst1wB+MTQs3lvqQA8YMUo6ZFMChGFcb
fwQestlbObmriEpmiuL183HmeeYdj8ZFpXDJHcRnMQFUvDViAldXifGrN+C0B930Nji3nhhfUHiB
aU09RrCu3JEb62Jb+6uItKX8/QKqjP6Ot/g2s8n2w0YfgbDC1kemq+D8BdXyJoX/JhH2/t4f4vaT
mr17iUvIojZ52/xFHSugOwnC9r0u033nD73/vXMhnLuJCm0XzjzISHN1xsImp7O1NSQznlrDjKD8
DvE+TEbszC2eKM8V48tlHi0J37HPr26kL2D9gQw2NIm1KZsPa2wLkrQvNIFki6IXg53TdQmeRYIN
EevkoX7hLzvVc5geqm4HnBILXHd7RRo9+v5+FbSS+5hK15fjgkPzWoCg/2AGRjbsmS7BpCeuwQ8n
EAwCiEV2atmXp2BXH7ySP9KYCOi7/WuO1K0bBCxFmCZYzVNXJcok3jhaAaOhVvbJruecJgWwieQd
09lGQmhxqW3us6pwodoTml0LcszAURoyCZZFNkEH2XzV8TBvnabEVTQ0qX/10zH97evz7jG69UNS
MBm+uv4evVmB6UFb7o/5Dn0ehlnmYvRgRoNJhJUqPWv7PKGmRsLLFzI1LmnwM2B74vnthIaRRyRs
RgcnSETrlbAdJyap47/E5VBXljAlWJafnzaYgs2OHj6TRKVQCrlebz1oM+61SbsgRDnDZAWl2sWt
Ri1IwMS2eKttdIrIJTYFm9prngQWnVYJ5ECcvZ2Tmt4rqERGBGt9lKYQa3P87pFr1DOsELjjnXx7
tEuJGh+oB/N0kTOjCLvxpv21QTF2Puvzu2w3VPkT1qrDrYlCJbu2oIBbkvngm40fE94HgEZERQkx
NsBP8Jy2R7lnM0pvAnHODw82rbWhU3A8dPWvuYxQDzPCKv6mRJB7R92RMqRIBB14iKn71pBnYSb7
j9vY3uGPO2wtfJmeU3uFYHY/+rFstonTJHG9voxCo2nyRRb1UNneCOOWrMgnZuwH91JaoD/dB410
xOoiSmuXTZ3JBJi2Lqx37vY1QXu2ik8bbJg7nTqsN2DFmquv2uVASfLm7BUJWXNx89uqGAVmmoN5
jc/tLSWilXpjn5FowBdk9j53RscJltI8pkJux+M67uAYfRYmfzt8l5DMPTVfcV+H26r2Wn+t8jz8
hAYj5+NM0l5ih1waqjUZGN0AnTc5i0VYKvzXaPkUI16KWnxJPjj8USvDscvgSRT8/VmVaJuI1tcn
k4auJeDmTwBBL5Qdsu3bR5zAsOgA086zCQYvuWfYz+8gTDSnyGRREQA2/mM+Mr8x1dNnWxdPVTcO
n8eXq3J00/nm+vvJE4QhKvYYwD07p6Um6Gyig6Abd0xR05n0WrTo48TsH7dt8t7uB67ke13r/XeY
s6PXxmLdc7Jhat6jP1aOBJ5dL/SYPVsFZu7zpagM2TooLHWd4PrQTa8IqszIuZgrnYiURD+Cuk5R
rrjcfi6XltNO511xkn/mNnja/jNr7lgL/Wzz51YXTyYXm1KYC3HhRG/1c9ApkFDWfq5rAIs1RdBV
gCOkEv/YRlkCLLlkc+Rbe9kZYYYV4WU5Ev9CFhCpv/npnk6hS9r+yUjQXbdvrBJ50pXsRisi81NK
E30BM6a4QwAV/rH8OhPMc+mOao7cycSo/JB927Mk+U3vWHROTpStAV1rQCkdNXei+w6LgY0UkdaQ
1YXELmpmKLVn7qjVOpA164BVXmSj8RXSpLmRBeqXB3rX+c1kee092tCTiTOm/XZsfUOedhwkKwWH
Tt8QnaLP+bL4bgVZM1R8O/iU6e6EIMllDcABokXt0r2W60vhZLILBtPkE0UK8Q3ikw6yfho48miA
qCXWljyzTGF1BOgkZ1WT9rJtlh6lNoXcYj8wxn3q/V1vPN9r9AnXGVkIVCLFpx9/AbogQGNcj+XR
y8hChkL5MTBaAM1LmVzBXanfsgX+lpShTv89a0TWSUnXrlkwIcNao7G//2uTAl3cWq5of0vNfWfS
znGgWgk0B57nY+OqVzGK12NVA1tvAmBEgNtWSeed/fpWws9brkgnyMy48J5unhxjUHstME9GbKoP
CNeAtvDY5W8pAffmnv4DlamZLhGL1gId4EC+5P1g6ngtHOTqWQjXSf1dO1GW1bKl9aw3vN34cJdX
TneAVBm0MKXFReo151eW2vU8suQldSX0/0bLSJ7IiEanaeILagaxFS+FqXgdZmtPjWPXzwUC8cSf
7b9uLFiotgJRGFnH/04y5hm0Z3mJ3QHVpXouMeuoy0F2JYLqRnUKklm4OhbOzLrxbdcJnJ+LvaSH
q+mfQ6sNtWJRA/689vpo5mv0pRkIjGKYAd0fihHkxBfC1NjjfB5QvWRCXqOj313REls7vcWzmwd9
+mHKvezdSdkpIVlDisXk1UJRsYb04tEc/xF2ebkuHxLRep8+xOHY16WXZMDjNnNWBx/NZ6CQlSda
Em28xlAJuD+WQ5xZRgS/oOqghclEfEt+r/CEnHazxQRJoVaGZv7YWZJxZS+uc3RaKO5Jwr5yGpNX
qLRy/GFxPSa+5l7MFe43FhrmjclhbYe+DIm4m/kKQiZPRBExHz+N/xVuhvpSW9Kii4CQTI/tPT1/
mTbzK5uFTh1bEPT+uEK/kpWoOaa/7RdcBFiQdTT+Lqomw52blWhhETKjjKJTSVCUXfXKUjTyproy
PREVg2EcO3stTDTWrDgrKX6Yw0/njCmJVNDpTLZ5WPdBSfJE0zg8jmAZ5VSLHVCwSu+wRRj++uw3
/HZXy6lyCfU1SEN6mUeJL+fImbIjUvvS2tMiIJ55cC8emorFBxMbbGDL0zHV9qBtmLYrug9tqGjG
O2Mk3mVJEZLAJpCaiSVMPDlcF9QrVM6wIkZsBgpoWh93hXyz+zWTeD30h8Vo2R/rxjUsuodmVr1t
QJadMtzOPKpH8Bf6y7B+Z4mXWzhDs+wRy2VqDCeqv/qJlaLzM+BL5ZrsUlhoSaOh8zlOr8BCO0Es
x/qegMGxl09fSg2LiO5OshqdPMMSaXS0XRuBjkgPcHDgDwidz4Q/FL6rCxgOmw/35MmPbhEJ5nQC
SJug/fbX5zel4QcE212KZj0/Mlg6Ll+ZepiW1LAn2J08gfB+opEpt4MjAvKErFESBgvSfd0KvjVX
D+SaDOu7LLAvAY7an7PxyVqKBjWYUume9VnwWzLdR9y3wps4e4n9IuJau4vBx8p5diLMRl7l9Nbm
GH5qJsvd29UgRCuyawMjNYeavl3CacG7cJzTIQeZWN8ic91BUDHWO8TYDVB/za7a6AiLbFskIhPS
KwQ8upxIWEUhwuEneYPhhy3US/fF/gZbONsjbopgIzrrxmQH/yZsDQsEISmLNGtVlSBtbRHYW5/x
7NoG5dh+6Wtmrb3RSDb445OZ4zCtvL1RR9mmSw1AISuLanVQz1NDR/hoUFw1VncHPU7Fk8xbm1jo
xfL/uJdzkKJ0ORUxlK4bljYIgVK/bwMWRDtdMGJByIun8P27NAIzU42TJ4n0FFgbVKZ6yyClw/1j
ZuunmYuaPisEPfC/N6ujWhY5vDSFACy4Dx8KW9WHivCGEQAjdlvzmyM6NXI+ukRqwnNUefgrvYMy
jcwl2CjiBytl8NJkK6ihSu7kScjkQxBX1IjpKkjSzuj829EzauaZG7jNByGTbUawphkgeztCAtdw
9caCJvvQOoYIZNYfchJ4NdZvcA5CtKiCmxj2mggggY3g+8u2FW/YNDsSa2RhaMRUaPjBuSOBhEYT
eeS4f8n+xpIDloLAWs2H04POul+kdfA+Zl5dIce8iOOP/TB5D0cOH6lTDY7EsGiP6X1RjfAKF1FI
prt6Sh/l5oMePoqQk6xhZaGyA7z+iJgYVIChdZRozVV4XByeO8skjEVcnv+XAaLeqZkKbS4FKs6f
Ns31cBcIJJNDL/XVHPLXnW0UubWdBxp94IJ7gtwc3l8anfd6ca8ysAnXygOJp28ATWKS+XxzpsUw
FIzqUPjIgM2JIgBtwI8trIaWPGkwh264aBwWSrCCVClPIGr7tduOcjfIqU81Z6oIzC0ruzISLxIJ
k9IVNyLWlldNhh93xtPKPL+LPCx+jeNilSguoyVe7XWDK3YhuS1oQy+Yx2Q63tAqfT4S6gv91BM7
Trqw+f/B05PphsB1rWYPrJbpSaqirfPDAn63ERbPwv5tEAl0YqzChoI3X5Eea7oMUwsXe8DmHdTM
cA+JtTEupxahCXwRbq3uWsSaThbNLw0hTxZrR9exszkOqywXdTy8pviUOXcavzmt7uJb+Z4UChju
ixTia6BJVX5aIepb5f3lTgwDt262jygmGgl29R0Y4mbVtH/25FKrrA4VHNT35WTlG/sSgJjQmlVO
dEVolaKGO/xlSMiaskCX1ki5UfcTx4feguf7R26a/1laCemJHRLdzs0QZMmGnIMD8iAcBnzEflNr
//xQqTAakS3izqfQVKXsASpOtwXCTyh0n4D//rXyyt3sujTc668YIW42VKPemq0Cft9iDCDe9Rp7
Ovj04BtEDHpPUnFRdZ8AFV15YJ7KNGOVoNBZBGswfA/TL+giSeslAyHLVDW7YFdU510AJEEKydDz
uztlg2Cs4zloD4fkWd2lgG3ey8ga3UdovGp0zgraJjUyUZiT3cFXSkzSgZVJat1zUVPFYaz3mbvc
SbCe6SHXfNsKhXMyZIOI0wPbuUPgTF8Q8tGwO2Ht2qQ8iaQueuOu7VrRvCBTMA5W7sAvBiOxyiSx
Qq6nJiKkDaVqvQypZgQgLuc7z6RFxpTwkBoT83HgvaJeRCekl7ZYzjxvywqprCBkU0nOVYLkTfhz
SGwR9c8n5/OCwDiUNtIhleEYFSlkAHhX+dB2XUx8bvt3LLLVVkrWE7I7Rf0C8zIEOPiKGQMmxRyh
BcZ9CFiPzbZjToLoENcFDgag+eqHgWUGA+Ah+dk7FrLJJUsFa1XyYLWtYp5XJmbJ04WyTG7D750a
UNVwFgkZTQxClpDDfJLXiGl0YmfDc8L0BD4ZKhAqStZuhCoYR9YR5qHOxJox0YpSRdaCuRbjCSSd
thQd59PX6LriDFjiwQ/sBHKjgYrvqaDphtZu8fvgKuji0lZ2xOYtV5B9M//sji04ThGy75liv1eJ
eXmVBGwBFYm875cPaM3AZDVHIenl/wKb8kIIvsmEn1HjZAAteN0EmNKcY7jfvLqnzFs0VtyxXzyp
0J5OUqlImrk5kO952g64hLH/f6wXUsdCMY5K8LxGpZCISI7YVhps4521pBbSbgZf4obQ1F5c6Vi2
oEcLSMRnNwsF+jx8ehzO5l+PKHL6eq44BEsPCm2LmjVBOu82XlZQlWdiUyiG0zYsbYNBUm/2gPMh
6JUpukt+GP+lSVJSLQCVHg+NECpzZ2nm+ixRM7hHger/LGaHYelyunZWyFd4iik7Cnz6lsoLDFnB
bqquXozbFYkuSnLuX9ZW1aACQDOW1Y0F1AdDDnfx0qSUzrDP4SrK1yvnZ+IsGd1llddkHhuHO9jt
KpolLhsTH5U0RNBH+iMy/+vlrHLJjOMKABq4vUVNX57uspJk12MUGrEI3aylwGL+qyUgG5EhxNwc
9p38ucGqnR1XQIXx0EHnywfrXinzhJARKZISiH6pFlsV6MRT6jxFH709l75hT6CdvmetdZK70PKH
npqLQ1OIPMA/AjqrcrP/4bQqkiSeLGbAC3UOLWeDfiLKIkSvRnO7yxL/62anUDwCfhuNVmAvd/Dz
Y80OodepqIyCzJEhHyrzuGR4klFde437G9ET2Dmr6gq+Y9LNlgkZvPFOQnc9i4JjLD0KV1nzIZLz
R/pPjwKh8AR16KNrT8nhO48p83gYonmsuRRSAU2NsSCA2VP1HPCwWgM2gr4At4/4kUifDzzl3rU8
SzOVc79wvFONcVxfEelloVdqguHbProYhUZA0Y2dXUTkKdNGjppweU0vbc1kTVg0O5G5cfyqxFHN
M5T9P5UaDrVWvqggscholLyPLKOyeF14chIdAerndsP+m0mwWI5gc7ZHCCQEYtYSgtVxotJ1f/jm
Nzeq9smGpJ/kHC2/BvRc5PYlam4ZG/zSsKFtsNlNnt9G/otcOAat/uwl+eArgvtnVMSziCI0oA/H
1xCctcnv/vfYlmkhnPrWZKI12UzSgKq6R4k8q3n/G3Ds/Xcv1+ETy2FAZGGUjhHOE3UjzifdyPjR
nSxUx2D7CXk+XmkHsKnQ9QaJvDP/4V5czsPU0UCHUDUMjnp5ToHfDsFBbdagF9IGJqO7GAdIGPYt
NjEyGpru6qn6UcfhBMmlNU7PbsUq8wBnocFKPEMTqBMuN5ni3ZKEz1hpiIU11SyoziKFXE/8pLXZ
f+OJ7ABKxLHfoa+qGpEqYlG+dpOasdfHcGB9XjsAt5Y2VeNCZ+Mrg0FdCrAvwK+4t3sdZqK8243z
xDz7NUC+IAaU98sJ6XFEHDRW3bgAN1PjdgWBApeMkLB7RRZTABjAuqTwwQ3wGf1bgehFLiloH5P1
1ouKG3hczzI4d1th77TvHrH3h7PvBR9e3lYkEPq/CxyOGXjRr6erOxN8kFVO37+fs6hSZ6RqLHfp
8Z05y3ihWNIFku+v9sN5sN9LZcKtBz+2P3NTTen4LoBERhFunpkDIeS0eTjvRjM1faAx894iQ7oM
7mayOsIzxC6PmkI6Nqt8aIt6QI5jpaiKdi+zz5NUS5ayICGh8Rul6br0+MqZ0ofyfYhRooRuTYMH
BF12JlH/DPlPLP595l+OqgjLxRjlVBojJlcRZ8kfT2baWUnHzXbwSz5/mIT5/g5klKSHPzSAqBty
BimonbdbgjrIedQr0tS/lHV4bM3I0N4xMxgI1JRtp4r4yPfVmqskarvs/r3QtrNPZ85BUF+AKpx0
nVletg1blug3PB+rl6KzJbLn4VdTzkU2zrW1pBnWYfQzxDs/9shLnLw+AQ4tIcZs8eSYRi22nHGT
n5q2byaPseNuivmCbRuowRf/rwyj6FAKbUtpFi2+mC/kWbOYaPALo9Y+uEMJy4ENddd61t4HFzJ5
6UddToBXbSwioqgfAL1nPjSuDsS8DSoaRkl5jRaL/dLqjBzyA4iMOkLhGCu+7uiBc8xpdVAXtPOI
3sdTMR08xd8iuQEE/BdhE14YCiPmmIH39hdfTFK8dya0uUEXtLPCFW6M/2fuCyHYYnR2xmLvuc+l
7MDlyJaUZ3gYGcRmLyWz6EpS96cnDqMg1RtKFj2Bq8213wylN7zDBYYsa3xwd1luwY2diHyZTz+k
WdqcMz67sDIhfUygvLno6glBvtvP13MEvxG0fuqhJyU81maFBdAuhjWs3LcuZgjydr2LHxJVeG44
kFKeICxG3UKvXdBd0KmnSYwr1elJWPyo+WtnPYKtzA9VWN9C77RFoIqhcIpynrUA8c5WtcfQTGol
9rRGZiV1KlAvEVH2XolKNSXf3vIp2r+QG3Y0T11Mi57az7V57u/jqDeXP6j9GuevWr7nUtKjpoTu
DPuYoZiDOumVPdqhoJ2lVVs6RN4bukw/a9+FG09V7iu/uUOMvFZFodJ7l2+W8fxBbdNeiqBtJY6N
xjVVHEUWeMBi/5lAr3JPLy7kTyKZgiK3e9BWx7k/Y1zV+vMM0U2nrcKM/qkl5p3EBeSGzROJUYwZ
THTaLglnx5eV9DvWuQUTT3soNRvZOTD1WthyypMwvBMhDTQ6V1PGu8iJTJBBwg7Q/5TtBoInSyps
n5bux5kCvxTIPcJr1qLQgg3XysdaGtiv7xi8fGz8aDEVlrY4a+Toi639m4034SD1ttAGsO/bkCnF
vIobQn61+eXVmxr8u/Qy/QbFR9SiJom7MdwzBXpC0ZF+8m8dWnTkz5HCveylkbH5dqUi9V54LNnl
1FyfwQgGplDfk0sy6/j09yfk2z8Up2vUe0HjR/CP1dWqXvpjcYRjHCm71zyi/XeP4xSAL4QR0o+4
tK4ypv8HVVvvzbsGczsaEruQfN+dGJBnn2mooFrKLqxh7bfsr13CKmAC2Pc0YuYuFMrx4jEq1K4u
Y+MeD6akxqVWikz6Df9f7TFJajaV/hDEh9fZfQoHSM6KSOfHB71u+2cpMUMvFLQBaW/Vo7NfPpyF
32htnBK1ZfjkfIOR7fD7aDiKAiH4HjSUly1pnZruDRNMW73TgWLwpV7E1iS0gCJ5XNi5Lng78gGf
CdBCs3TwrYoucDMLlAlWblv7ttY12T58nC+bWRPzc9sTg2PpmOMM/QKq9kZL9gwRVdpHFqEM+4Um
UYw4/Xuok00VNY0yDF8hSKj/veNuU2uuKBBhQtc0YLkw3mEM8ZZWn4YyMmxRDIePQn1R3zaM1k1z
LQdMz1TI0g/mTrEtNHsW03adfHxp7EMdM7nR/YwrWK1uO88iJ1EsX6sMnh3dpior6fMK1AGrlHD7
s7RLH3NQ5+yaH09QT6QLDK+oGPGGgO1ioFpyqr3lQN0fcS1vj7xq4ynEXDUEYdeEyf5+RPzsg+CE
BQNXAcT3Pz2MJXRuPpxRiK7H6jJsB2VyDCXsbqi9td5vZ7EwKknIV0sQB2Em3KBHHg1Oq3WGtcrF
gPcUX5OTm5JLQqsG0U3CWsLPKDYMRM/jupUJ9OoklTUR1a5WuGXVeTsrr2N3R/kbbY/anSm3kP/l
MzERsvZpgQZawnv/tjLRFeyirQWnwIlIKnlcSMoJaC9PShPAZMSj5gROcxPUX8LBahmxg1MmCfrv
Z9HFEJmtMhZBrpWCTYuq17BjJQTEqI8ssqdILx93BcpBAwMHtuhNObtsfQTIiFAATIn+tugmFTIL
sjICvjIwai1rxURNGxjwnNvTldApsAd1D3h5sWAIJ2MNlpjyktbTUAxNFEu1O1rHUfnTvpRChqnG
uymEkUZtAEKyrRY+iyySUPGcHg2URx13NKGV5VNBekYWdQU4WyYuywI3woiij1LnQ5R9MwA8Pv1t
JM7ugUQFGBjd/aU4T4XXobWEQp5RfqNxZz9CZ3WNcqD3/iU5nDLxl62ued6tJk3E53GqvNeNijGL
SeMLGftRanPdA6CTGlY1uwbvD+t1W595uNbGtNj7YhTcAdlI52g7syRql2xcNltw0mDKEPK41QsR
plWYoZ1MohKQ2XH4beu1oyS5RVGOAdyCCEoE0Imcjfknl5E3ktadc3JlAwIbVYZXQtJXSf73hgT2
Gl4kZ52G1g/3vQJT2YE+CggurUl07bhZEwXCbGOn52jS5dm+ohPtWz1o+wNzJvr1CbITyuGW1WoD
FRoIyP6+3+bZIueEN9kKf/GCKqmB+RSs9EmaUml61dddDlGMdjZpZXCz/A0qmrlv63JgJQaP2812
Uw/KdO6e5t6bYzbP1yqgKIbg6xLC6xDoFa2pENDorDo/PDSaatXthil/gxiPTMenk7HFt2cDInaB
PG80yxjkBMUGyMrROYA/+EuFUm5PjzeLaVqEuB9wKew0E33jjn0sRxC2yR9QQSQ5EG7Yel2gnWJB
cyNPhf6BCWUUSpAjr6O+aLifcjRYPeuS+F9IcpgtWrppqv5gWeZPIn516/xUu2Q8ez1FowmrH/m6
83oTfEBtYnl/bv0KhtsZnsSmObN/ebvEOnKh1KDBoFmb8Yz6qGyKfaIt8mi2KSWnmrZL63/0k34Z
tLCchCJ06V6aQNUtGMOp3xGqJhaEW7n5yO0PrRcpEEeChCzdrYkKXI1mv3yk62xcLpjrWU3M/+s3
iODOngGGtM6/MX/28ncaL2GHo+Znf8g9Lxoi3v6eAARE5D4xfQ47o5ELJv1jWFKHL8JFq70FO2mx
oGx5iV/csQHO+IJgJyw4mzdRII+hdLZ2egbs7xM+Iaw43vrP8T1mLRDufExJRteTafs8tVsfC7na
rkGc3IGao/g97EHuuSKmy06XyBBAFyzHLuLHPCPeudWrQfW2TWEyLWiXowsUa07MtEGoab7+vXNz
+MvO1uRbWKxOuHYxDmLrw3Yd4hS+66qWtIzXpfoVc7ifboSJxGti9ZemtYg4UzQ1IsUqTTzxQUZi
KflZ7myElic3WIwJn5Fsc1LkKjaAiWNbnEjIjBU/VAg3wzMgF0HRaot76Zm6S5pS94fBOWg9KUOm
1FhDoNBaNblqic/NIubSVsL8UMWHIzpM34NWfJAm5WNtlBHlezG22saB2EbqAg7jvXnMm6Mw02Ka
ap9FPS3G5uO7VNWHT+71loL2QhG5UZZP+JT0VgQdGWVK+hSgSlsq9G4zD/4w1T8pdt5dwjVUvVcP
degeNqnj69pSr5NW1SwFEmgjIQ1MXtrsIEm0RyLKIhi0fcbqisweoQ5imBfK8mGjRomFKLYW+nLm
jGY6nJMZawcy4OpvLWFHhpZLWtS8Hk0k6zYe1Yb5ufy/AqcmIYgHDKKsvSXOSeu8mLt8uaKIifsH
mDF2VfDE796N9xCyeAc5LieED05kTbTEFskZcrfpo65767IGF56D7QvzhWeZ4MrRGXd9a3jaj/yR
cRR1dn3z0bvtlrE2YPPWfIBh9mkJGVZe6EEA+9GE1ldYOryd/Nhn3wQy3H5wlGerlAFlg46LAmdp
ngLuxws3NSNBDv02SHH187UG/bVl3KOkV5xuhA3DDMsTgx7Sd6plLO5wD5zJsWTYEGR+ksY/dTwi
MFjgOeo4LDX3w6J2hoLpmexJnVubPlMYmAvl2El/oyefFCOl0BLFR2qJFcHovTAmu8xNqXekIKbp
Lcag3/2tn3iFHA5b86lNkrayn3fnhRyN8ak9lLBu2tGqU9h8UzoOdpACvKaI9qGkn2O5gWq/0vY/
U8QLY4cNWMTl5Ml+2w3jColXDJ08129PhcBP5FUffW+s+NOAkQeg1y9JDECifiIRMt1vAFxiPUVK
uMZQrZpfmv4qvhFc/uOlHByEpBznS28anaaljweFwXKpAx5sRuMPhK0IPAGibeI0f+APjIuv1qZ2
r9gLEo8peXHA2TDL/LWLpnMTL+w3wChunvbaLLskYj9MLocgI0wB5wo8W5pLZ/wfM8Xg1PhHhWm9
zeUXUX0ZbT5eR5s9w8ykSffpwqkCxWnBp2JJoLVtPYIcf0a0DAUk2nKMIZaCCmxbmv0p5cnVdE4N
N1WTXQPuh3AcyKSqfwuKM2F2kcKxPDTeQbk0V+iqnlG4nAM3msSvuxcw5ROHKUTv7bIAN0gtmobl
HBDY1bHxfoumDWpa5s6fh8vHJRT/vbkPi/z2kFy6G2aLg8IFAsLPqs44w9JokUPBlofipKuTlum3
f3HX9HuzYQsA4M1dpkNGZetokORWBSgPZSDEwVB/Vi7Q0c2kaYCU1YmU98oTerDALstWdPmpBaDg
VQ4cZ2asobj5OKtB2mXxx2hSQVhtAWpcuzBiH3dC+oL0FZ1qAV9rk479n3VYGrYKS3pSIcPvTnq2
si2M0DV/Pj607liZWXTRPNu5XT86v/JmrPpHfsLNS1TwMH7BYQkMCOQM64ZuteKYGEAIl+ZmzaZN
XzZYNb3VOshypXRLvtvvlkxHnOgipX0E1GmtXCqHR5cv/w+03uY/Gt4lJnOQ8DD/uab7N9pNmfuE
LSkqVg7ezEtQe+4KhJ+k0C9TScs4rAPQIH0EOhjANdWafTIStQ0BTN2fvm/Hw/grXz8e+EM7B+g9
28YU/U742Q6mXaO/82Wt5XWhUl0MFtZoHenIqVcidA91KxsOci/rxdNSVoF+Ma/ID8qQjtXNcSo7
Z521dPDsEG9t9MDUeQKBMU7+3R1F5T/8YTnuhtTMeKcs8yM2o8ys95OSLjhllUibHGGqmGHb1dKi
qcRUdmP6jcyGTWuAp8UDOnrKIRhZaJHGGhf/vcY4OFIeIC8Nd7Q3rO7s+23Dpk5tH+LGBXimjM8Z
I3ZxJ9snMla20unuwxOa3GeqkadpMPdz2LF/GiM76SKV+rldApv6mi453CLTNaojKjKykg7jdHWY
LurxC9W0OEy3med9bsHHoo9IWvhiIE5vhevPipulrqL5/BOofKeW6RfYXjEcPFPPap8B9uv+z0SE
A5vtLcKHVqD7P24QCga4NvadqWZyzvM4GW+YbVwGoGaZKoh3KFRox91BurtO/sC2zLk8yNmDWLEy
A3/A9oh5FjabL7t8J/eq/zvIc7VQ0fKp965cGE++MIIzDSr5P9SZpPS3BePMTa0XoRg3ZHSzcomg
Gl4OSsMJ+gQIAKnZmpdc1BpIolOwSdaqNwX2liKkx2PoXjFyGs4doZm4ro8RO7BCdeeYcdlvSHR8
V9lbtaVJDLhyr5t0V+8Q66fsSZvWdaYuIIouMXcTmO/2VPnWuATrbMTLvbHMAL4Xr18l9c07BFo2
Q/owjr5bzWrTofK5quGXTlqAiLmUfRFSfwjZUJYUZ+bRcLpZYTDQqHxvdcA7yuf6VvvuDt328itZ
AZbjZ0MbfbP5ilr8Tk/9ugYYCY24R9RqNchIrQSRhOAmmuz6PcWDTMKUuIyDc11kIu3XcNP4qohW
BOA+FblX/mgxaJHVJT1VyfLwHKWUa5Xuo4i3hFx/Q2OifvqqQKAsSjMcYjTT42ueB7NXDQJksYLO
+KSYfeg0K0kSIVUAIJIAfH+UDVvONmOSJeGPFSjndXGUYZBpIVXPwqwzhV4lx1vHp0VmvPgQDc2S
WUfG9GVBCgVVQWj1glCECOMdU+3w01qQWdOMmAD/HcyRR+7Y8d7EBKqBUNwMgd2I/zFOXUc0Gj8f
eRVuBr80ZsGHUu8808nQizl8mPCk/xPsN/M34QuksFInnzeBTdQ1ega2JHlTSH/AkBXrHebQ0CyY
ZlM9CrbJtM0R76VrC6YX8946UUBa6JJWSdAaoeHrLP3JtoHDGGd0+9CUq5uiENJVnp2QkVcSHQjg
mje95n3oEYY6UuuQa7zDqN77p95EY8kmIEFDFO9s2GEy5OSLdKwba6eeXX6C2Cw8gZqOV9ANEp+1
WHxi3IANWQ5nwI/9XHJn4ylWFAL85d2yA8AL6oDolr4pWKi7AS2OjanF0SGwE1k4cv+REPHPJW7G
JfzSeHsXU/llwO2/2KPe2fKo4hiP/sw0JGXofSYU1AX/uku+A8gW2g5lH8fTngKuj7uv2Y3RK2uo
IARFRcK0N05faHoij42jM2FqE38DXMhzSXS6lyHsd9HHVnRBJaichqJ6lduknhVbbAbZTIpAXgWb
HRUjUJn5dXz451NuvIF2zrfTwUWHJCygPkRZeDm2UzQ5mZl+9Y1KbZGy3Kjm8GZY5Tmn/ED8O1e/
G5L1OG/jQ3zGuGTSW4plfx+cAdJ1HU16wIxQTCRiSSU02qCuXthoGlFmrsd5TX8pVdnS1MdB2qru
6TE6wr5ESSNGkeZBdvEy8gSMNVAvb17yP5KbLhSJz5kAif2DH5oe+5w8kgcuT55aqjoNnhnlYkqI
Q+FstLb38cj189/7cbRVGBs1LSsj7lrzR/tTegfJbsLXAbLvtIyN/RcEgPmScVRJQJ66SIcyajrV
YmLnEiriCc9oQGNzs2HMkJCDdAlTmUdcUn8hYTBJA8eTILwTy7tpDpuUtEqaZ59SEKQLMU9zVSt1
Y46VmrHvUrdGWUcPww3lL0UBY2G79GuHOY67nS7DlfK3uH0jNucAkzLSvsLlFqXQqVq3SqdiCfUf
wJ1okqtuL+bmpFKw98nyfsWK0KAnMLzXAVhFtjfbHFGTlOK/BnvKZsp5FPgc3S/GjUaL/XxoAfvU
N341zW0+Zi/kck5vq/OZZlqnDOFJMwzaQIJaIlUFMo/nk1ks4rnIgtcUllCkFIjXUiMOkqNf6rzO
Eo/aTi2ofhiJcYihvvQL8Js9WVbWLhUfmYTkytfaryMerbAIj5RjQ/IExS2SKtK5SR3rn5npcQk2
2fPzPLqFpQFXZ1aNj8NGGfXjePiOmEN3kQ1rQT4M/H3AzXBipHa27FMPZQTobX6XKGelPQdeA/N7
Ucf34oT79YntabTX9hyMLUIMwhW0XYJMNyYGTyDOcK4DAbzD0IfLT+H7eLn7JwkN0lHgLUmuLtDp
xEjcTyl7O/U+RQzxO0EVmDeKw0NLUV1TRWDoW0rB8rGecFLq0jaQOMQXK/fWW7TduyKBzVnyOcrs
Urv40LxKYOVzlR4Gkl4RfSKoDzEkPg+GosflIrC+s1zXHvsu8ZC5d87WCfPrYmlO8ffgK0RipPtD
xIt64CYerJ1di5B4RSodFWTCfIX1j7V767+PzLaBlkl/S/8aeNefx+B/LUID1hUuRmcHkKIW/Dur
9TbdZXQTQ8qdNTqbzjF46m1W083AYox/+Y1kH4udP2KkIdbQPyPYCSeJHC6OrArQsa92GROsax97
ldku+AMBLvHQPh1NAUYIRMStiTgk66J01MJNCjS7d7pTdno9EtS+l30J9C1HMI/u26gX0m1Okvdj
avmukAmXy0cOjUJHyYM+lTpufzPAyXjg+84zBuXnpa/DDjPT2bCig6fYdl+t4SQeNdLZxmG0FCmJ
4p4gO1BYsQRPmL3gfiRNFqfWLJGA7GSI6bemO7HTIcVtGCFTARUjLgz92n/ANRcIG0DOgOoDCS6R
MsY7vNURO2SbRF0r8TGs/lF0/djFoIZFqN6TJuMb0YluaamWKcKj9sNOoDz1w62EP/+TWB/AFgxt
d5vJsbd/nEBLejlZ7cA5JxmvThpz60v6mVHvLndTJ/3FdUqvPSZviyw1vM4PjnRuQNcc1VZc5fM4
9KO2yfTObaM19qOS6zdVHDu1VsycXWRYFX6pm2ZT0vZIHOdqn99R+pVqNJWyJRIvKnAhEg/HA7hG
Gzhj4+yfrmoy62lqdG+cTHQqh5qbZjkGxMNvbLeX2appwHZBq2vh1wmFUiwrjc7cLgF+ZOx81RSN
D3b3zOipAfpl+Oj7/lgg5NEVN1je2GMlR4zqy9JslcBPiTq3H5aWHUqr7SQvcFv3mbG0EhLqJwuH
j9VjyPb2JCKQipfKUd4mddQLb1s2e0QQ9ujNcug1gnxwT2w6nlmu/3Ty+lq+CaVqsaV/sqppmzln
VNuGOgbkL38nqSWJW9yCqf2Y9XmZKKd55AFQJ9Fwbzz1stK3C5uXgza1Cfurp2lK+pJ8ci2J9bz9
mUwTindsmuupxwNdTEVYtUPq9h53sq1v1CXcExC4RDvS8CLYKzsNi/sFuI0iD98lMzu2qe61fQYl
gypEjb8pFRWtheh9qOpEO+n+Z6attUiphyQupv6YplfGv67JSN/Jtz15udHLXkinjuS+f46WiQID
MWNk9/Ftn5pxlhflNptFMRkbpzJ9fdGgJbLj9pGtVE+2v8Npu+cLWEd2gYD0S9ipgWOWhTyMzrAq
BeCFF666J67t0XWaud6fkMIOn4F7WCBqoZE7umCMOxDBN1PZERclgq5YVM121RHnDz6aY+6/gh1g
8fLIRMgy8NEFzzCaJb9D5yNgSRbJoZdfXYubJaUHWHqhTredXGcdZvPiTZ5653P4V3wyjQEl9/kg
SRoiePZ7OxTK9RXsbRAvFn+sO94gKW5MeyGb4lIORxU/+AzEC+/J7y2EzhUICfX4nl+A6K2v7LoF
3OOIFkKd9W96tjicgI5L4W7M+84otICp/P9KgrSGQh4/6biJT5vZprvR4JzIWwnEei7cvwg8C9OC
uxmbMga0BIfgtZ9OPkYwxVOEMxGtmf3m+WT0/+pTrRtzUckyF5xkncv+Cxyn/b7PrQ23u+Y5amzM
K4xUW25jPUMBwyGBtNzYhUihKtpkGIKODfBfxt6aZeOwccQ/LN8iyuMgUgMIycLP9Fs++LFH6Kbz
A7jiDcTk3tSddq8kTMz/Hp6Ffv8yB0B3U1jOAorzDUz85Gy+I1XE2iryulyTztzCeMoFfXwq2J0o
3gGyhCgfuwgpXhzrz2UM5iFLGaQglcu6bMhOavz826rB6nF9+jbBVfJuekzsGq6VV4i3MXNVYPFm
AEtsNdSBiJ9Zig7YxG4C5T8c5Kg5THwy26vSERdPInwIordF18mrlqNyXAn523LaxVn8kbVEl8S1
lR48/6aLY0wJNEGImR6R1USV3CvXM2fy7uPrJoEj9yxCC5fytDuc8JXuJSWrTpbQ0ItLAuh+5cgU
yKqC4AGy/ayMJi7E4BhqECoh1ZMiNcqxTBtQ9+8o4WnDOLw0PHicxQkbtHrYeiJQhsQz2lOzy7kZ
FZTInmrJfewPX088ZJok7jJ/KDADkFxR9IlcoDi81YcB39Moy99358B1Bq+W+DL9g2ZdcI68FBCP
dJDKuFfGr2Kf8E6IgdmT4aM6dHZga7u0xOhGpT9OfSMcWwdJ8UB6g8PS/ypisCXgbSCQ4a7/Etna
KhlYACJmcBd1bQTwcWhaagTnZ/Y4U+8iGb18cOQeyp7peXKLyQWFEpWa8hzwVIYUwx/re6BAz6Cm
Cbyh0zR5u74YKcRfzc4mmpcx1AYyFJOCYuoGdm6F15rBFUcfuwZ8uzYYQRzp10umQ8YFkQ9EB385
SOnG9/D4Eh48WlW3ik/dDCVV3JdxLw3pd60sgjD/oTPzbQmI0jti8wHYx2CV2AUZCG75gom8WWVW
u88XMIEcw3ptAl3JkSVXGl9p/G+KAM9c4jPUd7NyWCAgSQoK034IIQM3x9n3ecQDW/SNcgZP9Bbq
BRocdcQP4tN8I5XBfqAlc7wMAT0QH9gBbBb000s/ypag6OxqB4dWuVI5l3JQdyi69p9YvscJW4GM
NpScRIBX5Wsb4Hami28pzP4XNJFxjYKMT8/ty0/5NFy4zRwDeTmLfjy2tIo4y8MYf3I300asQnty
6kU1VHPeDChHG3a1nLiOVQ2gePPBPBh3FhPCcWs76YThp6XHJaGS4UcQC3MdoFCC9jsNb0etwnr7
NE4AgYhGLWWDa893HjglX3vl4C35aLETfAkpXCr/UDfbKi61DN0i4DL4n7aCKg7DNqZgRbFzISGT
FPCXNxXb60uVJcx62xJcrR2Hf/yeSy1iASQeeJlEHyGN4HJ6yZaYeotVPfdEedgnFvFN9TnBGZQQ
JqK0qGmx7yiX8/BEkVkxbaVWoyVHzE4MNslGOMR4cO0N7vwc/PpykpcsWPPVKLjEqJvvAjBMaHrq
Y4m2B3AWAJROwWB5Ar4IEu1AmuyXo16uDjdX/ZYWg98JgP3pgFnOW5Si88CBAwXIW+Ca9e4xT66Y
FGVTgsa278mTBBy0P58jOROZIjovp2ipNPQEXJYzyVa4P/CVv0Xm6LD0wDWMrjTlJxx0JO0OHSHU
GFCZmDU7sWeszuDNHPqS3EGqQhAPaett9skYZ8PEOnG0bOuYiMjYwFVMwgLHqp+QPZU014F4fkSu
Ezm5pD2WbYGye6Ftu6+Y14e4qSjuIoZ6+r7lDwGJzEpYGp7cuM3pQzRgz91LOzUILneqpAubU9zV
lj3a5hQbnF7lIfooScevvnW3e2ZiIHwz9c1wgNjEI0nOf+5b9GEzyN7mOZKhDxzKSjBn2aGBXZYw
YTcc36Oe3Xgu+MiO5EiWvZ4p4oDnaYylQpmNUlbl/AN5uhTJTBwruxzLp8OCXKKoOfoI44xdf2ct
WaIZWrlmDfuQvpgq7bvzeLh5f/6nhd65uZqTMHUbm279cxwG9mWBbwrzMtCShG8uX+pAZrFGfpFo
zYOs/6iY0pg6S3p0HzXsgl1rFyDv+a7nlgYU0WJnfnKncatXM5v1jkcMtznHG0ktK5AA/vD1s/Ap
wXYqfZD6SF+VFgoi1JTEuSOtP02UFN/zOSXhnJGWL37KH0Mmpn/3FDatuvi8CDIwsnn1em5DAIwM
mqVLjqka9M6etbp5ftvXLDgTIjkRgj+4UOc5FdBvho83USOO86S5/yivAJLfCJdiRPZepCrJqBOW
PDALhLFqWSQb1+XTU+OHCJZlH47Xv/g4ISdAZImkmN0nP2rg76kN6M3CQEQddFvO3gTY5NjWVY3J
jZwgnLmScozR8wjINDst1gk8F7Z2v4AmeTf4UuDFgMpyMcS1rRF54UYv8m3x6AcsR7ZASABwtE03
p5TqjKenM32US/11lEKG/+maDGDUvoAQFXNbv8WZwHnMGM9PywthBURmgHBPpqSABAEIk7GR0LZl
MNraVEt2hwRM3sZ46q/TrdIpc88yN59uchZyw511pJWBTU+c+4zIwnj0dAkW39zQsKWhSChIwrUu
EJqnaibuqfNUmLwar7kRJVdBLtWTd0lUD0s2aqhP7o15qM7MR1SAsAauInTE0NWvFfFeV93AE3Ta
WPXEIRuyISMIdeOzZKsuMJTdYsaALyLPWaJs+8bsgLFlhRga2ZjEfEtogNXQLr8ttx/Qn86kcJR8
fZC4UemgsrlqncevDOMDBwX96OVaVlkSOnWg3fFMHZPstcG1sS11e9XtUWUacVBd6674gd6qb5eU
cbBdb2Su3qwEQFwa9uJumjEV+eDJX0JIGLGjazU/UNLvzdPVyT/829DQAWEtrUrXCbDcY3Q9xOa0
g+YhlkS712ljm7bYbgRrk9S4plIbInDeyKmCX0MQDPvpeigu1dWNeyu2d8PmlNhuiSLiRkNQbTTg
L85KMe4303FT0uOnI8S7gsOy8XLhJj2RaH2LDTV35uVtmb0n0UAYqJQlrmXmAxXP1bN9NXo+qBcc
bIgIsJlN6OqinV9JSeOt9e9SWX9//QqHEasg8UgI5Dgv5ret3ma+s5woupBXcjhldsq+zv33IriY
Q7rAbMpcwnJkZLdneDABfKOai9tRUAVX13Ttd+IjMvDnV86HRcM9TZiR4qHc7dKirFyW5ghL5f60
+5BKzN+I4dQLDCJjOz6b2OPSA0Wsmm9j+NooKFElesWBgPhS+55c//y99gh2uCWcWHrz1p4S0dwc
qAEut7jV9SH3AVkXDj3yeaZb8NDrCEkO3KYrFxEDa+sn3Gr54wipb0KXtu8FItHfg2v6PmJk0Eo7
VeIEuYtJ8YUQGJvRoP7kU5zqVKcKa56/PUXu5Zifsyw5CIQSXjuMQIw1vna+uaR01pIdZCC8UCbO
snXE/usRvFT34wqBfIbh3lkOEQmH0pMS6/Ro8WUXXMulUA5mdqbaa8DbxwQU3q+dUUjKn1Clk7OS
tVyNw8eGr6v8VXU7ENcJZZoaMJ6sh+rkr73iZVYzhm4blb23pmAs3YuAEd36JfrNguiu3gCd9BZM
XoxAT58Q8YjbLHTtXDSr9gUg9J37KVOGSe4z9EfDpkGkvLcdOa9iHEgphGpMGUuCmmv0ZyEcBgTa
Zb4S/RbMeZnqlT6i8jN15IbZR2hrZBnQIqHlNLcoOrwkm8rVgNS+c6N7RgpBnGcB21n+eUtFX4vY
7U/7ugi3EjsfxtXAcPh3/zr0d/zLXYhRBagrxrFCDuvGmCOHBiQREdH8H86bovby+H46xxAdrGSd
9d9LrFb0ASjrPwaTf3YQGo8/4KTcNkd6JizaZ4S7iGO7isCv+Kkm59CkQHjGQ4e5OqxdL8fEmsYj
YbmnoaTNRyhrY2ug2FdG9KA0bk8ENShMXPiIHX+B8+OVgoj52c3Y+sAggrptTYqUo776SQWjBr7+
XtwauvE96MOYC/LPTE29/t+w9tzM680/5vmrQY6CG/+vuja9+0OOR8RX6psCTcLJQSZzPGHP60s7
K5rW1mM/9xqpCgMz1FNsGhsKTxJw4MExUeDR7eHep2GrWzKUty00pPuj/sQj3+FnYjejU/U2sMmi
wS7UIt0P9+qbz+veQG6n0pkreJGIc36/nv+hQUZ7gfcXVf5GZkYtdK4WEsiNPDf9snIliz9WOLYB
SjbC6NVKbnvJbbX6hNCcCHpgC+7Jc2zHefvOd8U4nkQXknFfvMpo9+qWGsha0c7Aq1nZg82Swwqn
Kbum0rfBQSQvo/3UeWf7OcomBvNX/x9FJ0BuH0A0ODwqIx4fsYoMTnZeIkOIQ1rXhbbu7oc4A9ro
D+2am/2Ub9j/gz0A1ijgY7CYcLOrKJV+vH4i2VYXLqz4FUDnwljDJOiFYR8ZlDrZ+mnmfibG9XLO
9KkViFQMfzCjzEknaNTKdP/Po7SAlnJZg3KkkoVL9/f6LIqp3g8DXrojFrO3KlTjsAWFTKQZrMbI
E7zKA9u6IUf8smoKr80fewillkAU7vH8OT4l3+lYdhssGsjM7N1FNo8q/QqNzX0ofMbUEJiBL3xF
41nJznziGqLVRaTbAbaZAUyt1gMN9FA0bpTawEd3zDibsYGMAhDdypOosIctcBQGQEllGkh11PeT
3jnhpr9CIFlNck/BpenEcm7m8rBfwvb3qX/zTDxLN9NmN4Jqn5skYnx2Y0+BRMMzUtE9IfoROXKc
P5jab7Q6g9w/xviGqpP0jsfIy2cXNifbb1i/b9TCuqJ5qd0FrmAF6Crz8xnJwU0go3SHAK7v9p4j
5P+QrU7anki3piTEXLbJNqO8uT44ioPjtI48d3FMYjjpUar9L6S/oUm6KX9pVuMrKH3um2hPDbMO
Uy1AlCAvdQJKjoJVmoROv9x5pnEbECvTc63W30m0mWOOtaQ1LzzKjQrfTHff8NEBg9EsxlnZ6OTs
xtYLiKowlbgZ6aLQfi7I5airtdmBvKAbjJr8c+aDpBBgc4L9gx8m7HcX8GUKLN63IoE8H9a+kwJz
x+0+aN2Yrx48erpFbwk9xbDOA1Ih9377hHHvdOQcH/ZcB+uXsONgYYodOgyzOfh2Q26xaAy1+pXM
pWJwpVbKqOk5SLRQrtkVrHxRSmaQp5qH3rvZezbhVA47I7XrcObEmT2oftRe/KQU686jqXIWOBrY
ISpw+jypCaJek9eDJ6m0bdeeIJXqHnLA/rPCITYCHw6jkW8OFD6TKnxmIFLXNVgUf0QTCTwtw9vz
MfRPthz4aVM/JyYSJpxEz9qHZrbQAflWlAJm5BOKLk9kj2wR67Jf3fzpHxnD6FCU3JUB+MzbwnBM
MrPs6ScqcRZuzEKG7oQKSvMDRAyjjcC7lHalfVJ5fmgJzSqrQZ3Mm3j2OcM7TkAZKvKUrIjEBOkv
ScsytnvU8NEE7phOXeQ+HDNKvEeA43UgWCEAj2oqAX3G9ApJhUs/sEnZv6BJFed4jqNulnLk4MrX
Abq7an94YompqjT4S5n6KfbikYkJiCHx4yVpfkIgf4RyhQwkXUkjIRWktqp8hTR1zlUOGGab5wd0
E7pYC5p5hWHdBUFg7SIxuTJnIUaWBnpUwQGPPThr4DYKlzkkPz9GyFQlnswda6qDdeASUW/frvKg
AHuImxTHKJAXf+mr3TKMrjXv7BdNeIo7DQO+VfdjOxg0WwRls/6GguNMyCmqEwfrlYJvL9doizpw
p5Yi0PhjG9k956rEYQzuhE+cH5WW2s2HM24t2NxBIsoTHs2UAx8wnIrkI/mEomNIphWekX22//h4
m3TJIbxtNd0XJg+vgMABELlIAutCi5+hsgZmi737PRGKlAugiwWptwFg8g2T5Q3KSbwyhptKej+F
FqnuS+jBe40RCZ0Al3xI0KUOzzJHaNa6n23cVcIKYE0Bjrvkn8SqV2Xn3jz5OqTtTN2bx/8ZjFgb
bk4XL+/dyvsVQseAzDDs5Uf97dOe0LAEKMB3+NTUQjLIpQhKiA0dopZSL4TW48BkljhY8Rdr+V5c
BDli52S9r9T6+Q2HQrkC6CZBW+SswhErE9vU5+PRZN5zrWGskFiQ7QgMNt5aXA8MjVMU/SW9+Hf2
OQEOYAbIF62/4fkmyC+PGe+LY+lU8uN3zBpsCZKNRVRIySLeE99c6rxekb6q5nDNL9aOmifp6yNV
eJObtHXg0rlUof0RJGjSQLCd/MZ35eQH95KXdzk8qOopZyWNMaEtZkzynZ7skf3UHvJu+8btgeth
77riXQ1ThXeuV9pKwG1CNxaGPt9YTEaNd7VufUHE4o4z6Y2AeasUzNuXAeS1GIcqRR3e3NC5yYbO
Hl7dlJC1m8XmNb/BzM+SnE0PHJYoaP+0A6YmHx1OjFp1AwfHEin8BIPlMDv3cm+sqKkvKTC3umQd
kd4zYJV/XdX/jAzFSu24x/MjVjFF8P7zBOn88iR39Rno2DxAyxZPfvn+JZjeGOzUMAof35c4DNiK
03wgjiH4TQMAWL3sgHxFt97BOHyehGfNUC1uxl6lv/aTkGH+B3vNzSoCWyHEiypzbe/knkm1z1oV
bltsVueRP2oNleZY5/EN8t8UUZSs9Ou7pcgg+nkAv9cB+pY55s3LfcY5pdyZp6EoWb+7HNJZJMpb
upb/mzZ6oZnveTXf/pG0qHdjCBuYBB7O7siC40XGh+hKGGkevX14TxF77A9mxYK7Ifk1llSn9Wmb
DwRttkqNyh9KrtJYq14Dt+vRr7cdrR7MyQlgkB63mFO9vNsGbyNhAV89lyQeKkkxecIOzw2IP95w
iJn8HstlzJQmTT8J8tx5JDxJFgpnxgC9YDQsZQdisbSp6KnqjKwRyK1bCyiDadZNOppcw7DhFU3v
9zbgrGLPU6VZFtAISRZC+L8UpItelfqtIcEq6cNi5uaD5gzsneqo2nvCTwhkoID6MzZ8Li3O8YQ+
VNcYDsKpK9luWu0vVZ70W6HkjhaRZlaO3JKhpU6KexP7O7jOSpx/8A4L1xD4Lx/DJNpNUGHfdyuk
m3FZQIRFZCuJjkdZN6EoHwIqsEwEpNkRrEANs3dL4BytxjQcwUUtyVQUjs37Ty73e/00tNuftCQ6
oU0shFzDWKfWcNwD1tYXoxrwuX8fFpQzNDVRavSy7egm7vRS8YgXFM0IVsvluCMgDDHb/9TAXQYy
teOgNdaRWsw8+0T6iv3qTt9xtK1ide3qpqo=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw5a;
use gw5a.components.all;

entity FP_Mult_Top is
port(
  clk :  in std_logic;
  rstn :  in std_logic;
  data_a :  in std_logic_vector(31 downto 0);
  data_b :  in std_logic_vector(31 downto 0);
  result :  out std_logic_vector(31 downto 0));
end FP_Mult_Top;
architecture beh of FP_Mult_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \(FP_Mult)/(FP_Mult_Top)\
port(
  clk: in std_logic;
  VCC_0: in std_logic;
  GND_0: in std_logic;
  rstn: in std_logic;
  data_b : in std_logic_vector(31 downto 0);
  data_a : in std_logic_vector(31 downto 0);
  result : out std_logic_vector(31 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_2: GSR
port map (
  GSRI => VCC_0);
FP_Mult_inst: \(FP_Mult)/(FP_Mult_Top)\
port map(
  clk => clk,
  VCC_0 => VCC_0,
  GND_0 => GND_0,
  rstn => rstn,
  data_b(31 downto 0) => data_b(31 downto 0),
  data_a(31 downto 0) => data_a(31 downto 0),
  result(31 downto 0) => result(31 downto 0));
end beh;
