`define MODULE_NAME FP_Add_Sub_Top
`define ADD_SUB
`define NO_CE
